module sber_logo_rom (
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(128 * 128)];

  assign word = rom[addr];

  initial begin
    $readmemh ("../../figures/coe/sber_logo.hex",rom);
    /*
    rom[0    ] = 12'h000;
    rom[1    ] = 12'h000;
    rom[2    ] = 12'h000;
    rom[3    ] = 12'h000;
    rom[4    ] = 12'h000;
    rom[5    ] = 12'h000;
    rom[6    ] = 12'h000;
    rom[7    ] = 12'h000;
    rom[8    ] = 12'h000;
    rom[9    ] = 12'h000;
    rom[10   ] = 12'h000;
    rom[11   ] = 12'h000;
    rom[12   ] = 12'h000;
    rom[13   ] = 12'h000;
    rom[14   ] = 12'h000;
    rom[15   ] = 12'h000;
    rom[16   ] = 12'h000;
    rom[17   ] = 12'h000;
    rom[18   ] = 12'h000;
    rom[19   ] = 12'h000;
    rom[20   ] = 12'h000;
    rom[21   ] = 12'h000;
    rom[22   ] = 12'h000;
    rom[23   ] = 12'h000;
    rom[24   ] = 12'h000;
    rom[25   ] = 12'h000;
    rom[26   ] = 12'h000;
    rom[27   ] = 12'h000;
    rom[28   ] = 12'h000;
    rom[29   ] = 12'h000;
    rom[30   ] = 12'h000;
    rom[31   ] = 12'h000;
    rom[32   ] = 12'h000;
    rom[33   ] = 12'h000;
    rom[34   ] = 12'h000;
    rom[35   ] = 12'h000;
    rom[36   ] = 12'h000;
    rom[37   ] = 12'h000;
    rom[38   ] = 12'h000;
    rom[39   ] = 12'h000;
    rom[40   ] = 12'h000;
    rom[41   ] = 12'h000;
    rom[42   ] = 12'h000;
    rom[43   ] = 12'h000;
    rom[44   ] = 12'h000;
    rom[45   ] = 12'h000;
    rom[46   ] = 12'h000;
    rom[47   ] = 12'h000;
    rom[48   ] = 12'h000;
    rom[49   ] = 12'h000;
    rom[50   ] = 12'h000;
    rom[51   ] = 12'h000;
    rom[52   ] = 12'h000;
    rom[53   ] = 12'h000;
    rom[54   ] = 12'h000;
    rom[55   ] = 12'h000;
    rom[56   ] = 12'h000;
    rom[57   ] = 12'he90;
    rom[58   ] = 12'he90;
    rom[59   ] = 12'he90;
    rom[60   ] = 12'he90;
    rom[61   ] = 12'he90;
    rom[62   ] = 12'he90;
    rom[63   ] = 12'he90;
    rom[64   ] = 12'he90;
    rom[65   ] = 12'he90;
    rom[66   ] = 12'he90;
    rom[67   ] = 12'he90;
    rom[68   ] = 12'he90;
    rom[69   ] = 12'he90;
    rom[70   ] = 12'he90;
    rom[71   ] = 12'he90;
    rom[72   ] = 12'h000;
    rom[73   ] = 12'h000;
    rom[74   ] = 12'h000;
    rom[75   ] = 12'h000;
    rom[76   ] = 12'h000;
    rom[77   ] = 12'h000;
    rom[78   ] = 12'h000;
    rom[79   ] = 12'h000;
    rom[80   ] = 12'h000;
    rom[81   ] = 12'h000;
    rom[82   ] = 12'h000;
    rom[83   ] = 12'h000;
    rom[84   ] = 12'h000;
    rom[85   ] = 12'h000;
    rom[86   ] = 12'h000;
    rom[87   ] = 12'h000;
    rom[88   ] = 12'h000;
    rom[89   ] = 12'h000;
    rom[90   ] = 12'h000;
    rom[91   ] = 12'h000;
    rom[92   ] = 12'h000;
    rom[93   ] = 12'h000;
    rom[94   ] = 12'h000;
    rom[95   ] = 12'h000;
    rom[96   ] = 12'h000;
    rom[97   ] = 12'h000;
    rom[98   ] = 12'h000;
    rom[99   ] = 12'h000;
    rom[100  ] = 12'h000;
    rom[101  ] = 12'h000;
    rom[102  ] = 12'h000;
    rom[103  ] = 12'h000;
    rom[104  ] = 12'h000;
    rom[105  ] = 12'h000;
    rom[106  ] = 12'h000;
    rom[107  ] = 12'h000;
    rom[108  ] = 12'h000;
    rom[109  ] = 12'h000;
    rom[110  ] = 12'h000;
    rom[111  ] = 12'h000;
    rom[112  ] = 12'h000;
    rom[113  ] = 12'h000;
    rom[114  ] = 12'h000;
    rom[115  ] = 12'h000;
    rom[116  ] = 12'h000;
    rom[117  ] = 12'h000;
    rom[118  ] = 12'h000;
    rom[119  ] = 12'h000;
    rom[120  ] = 12'h000;
    rom[121  ] = 12'h000;
    rom[122  ] = 12'h000;
    rom[123  ] = 12'h000;
    rom[124  ] = 12'h000;
    rom[125  ] = 12'h000;
    rom[126  ] = 12'h000;
    rom[127  ] = 12'h000;
    rom[128  ] = 12'h000;
    rom[129  ] = 12'h000;
    rom[130  ] = 12'h000;
    rom[131  ] = 12'h000;
    rom[132  ] = 12'h000;
    rom[133  ] = 12'h000;
    rom[134  ] = 12'h000;
    rom[135  ] = 12'h000;
    rom[136  ] = 12'h000;
    rom[137  ] = 12'h000;
    rom[138  ] = 12'h000;
    rom[139  ] = 12'h000;
    rom[140  ] = 12'h000;
    rom[141  ] = 12'h000;
    rom[142  ] = 12'h000;
    rom[143  ] = 12'h000;
    rom[144  ] = 12'h000;
    rom[145  ] = 12'h000;
    rom[146  ] = 12'h000;
    rom[147  ] = 12'h000;
    rom[148  ] = 12'h000;
    rom[149  ] = 12'h000;
    rom[150  ] = 12'h000;
    rom[151  ] = 12'h000;
    rom[152  ] = 12'h000;
    rom[153  ] = 12'h000;
    rom[154  ] = 12'h000;
    rom[155  ] = 12'h000;
    rom[156  ] = 12'h000;
    rom[157  ] = 12'h000;
    rom[158  ] = 12'h000;
    rom[159  ] = 12'h000;
    rom[160  ] = 12'h000;
    rom[161  ] = 12'h000;
    rom[162  ] = 12'h000;
    rom[163  ] = 12'h000;
    rom[164  ] = 12'h000;
    rom[165  ] = 12'h000;
    rom[166  ] = 12'h000;
    rom[167  ] = 12'h000;
    rom[168  ] = 12'h000;
    rom[169  ] = 12'h000;
    rom[170  ] = 12'h000;
    rom[171  ] = 12'h000;
    rom[172  ] = 12'h000;
    rom[173  ] = 12'h000;
    rom[174  ] = 12'h000;
    rom[175  ] = 12'h000;
    rom[176  ] = 12'h000;
    rom[177  ] = 12'h000;
    rom[178  ] = 12'h000;
    rom[179  ] = 12'hf90;
    rom[180  ] = 12'he90;
    rom[181  ] = 12'he90;
    rom[182  ] = 12'he90;
    rom[183  ] = 12'he90;
    rom[184  ] = 12'he90;
    rom[185  ] = 12'he90;
    rom[186  ] = 12'he90;
    rom[187  ] = 12'he90;
    rom[188  ] = 12'he90;
    rom[189  ] = 12'he90;
    rom[190  ] = 12'he90;
    rom[191  ] = 12'he90;
    rom[192  ] = 12'he90;
    rom[193  ] = 12'he90;
    rom[194  ] = 12'he90;
    rom[195  ] = 12'he90;
    rom[196  ] = 12'he90;
    rom[197  ] = 12'he90;
    rom[198  ] = 12'he90;
    rom[199  ] = 12'he90;
    rom[200  ] = 12'he80;
    rom[201  ] = 12'he80;
    rom[202  ] = 12'he80;
    rom[203  ] = 12'he80;
    rom[204  ] = 12'he80;
    rom[205  ] = 12'hd80;
    rom[206  ] = 12'h000;
    rom[207  ] = 12'h000;
    rom[208  ] = 12'h000;
    rom[209  ] = 12'h000;
    rom[210  ] = 12'h000;
    rom[211  ] = 12'h000;
    rom[212  ] = 12'h000;
    rom[213  ] = 12'h000;
    rom[214  ] = 12'h000;
    rom[215  ] = 12'h000;
    rom[216  ] = 12'h000;
    rom[217  ] = 12'h000;
    rom[218  ] = 12'h000;
    rom[219  ] = 12'h000;
    rom[220  ] = 12'h000;
    rom[221  ] = 12'h000;
    rom[222  ] = 12'h000;
    rom[223  ] = 12'h000;
    rom[224  ] = 12'h000;
    rom[225  ] = 12'h000;
    rom[226  ] = 12'h000;
    rom[227  ] = 12'h000;
    rom[228  ] = 12'h000;
    rom[229  ] = 12'h000;
    rom[230  ] = 12'h000;
    rom[231  ] = 12'h000;
    rom[232  ] = 12'h000;
    rom[233  ] = 12'h000;
    rom[234  ] = 12'h000;
    rom[235  ] = 12'h000;
    rom[236  ] = 12'h000;
    rom[237  ] = 12'h000;
    rom[238  ] = 12'h000;
    rom[239  ] = 12'h000;
    rom[240  ] = 12'h000;
    rom[241  ] = 12'h000;
    rom[242  ] = 12'h000;
    rom[243  ] = 12'h000;
    rom[244  ] = 12'h000;
    rom[245  ] = 12'h000;
    rom[246  ] = 12'h000;
    rom[247  ] = 12'h000;
    rom[248  ] = 12'h000;
    rom[249  ] = 12'h000;
    rom[250  ] = 12'h000;
    rom[251  ] = 12'h000;
    rom[252  ] = 12'h000;
    rom[253  ] = 12'h000;
    rom[254  ] = 12'h000;
    rom[255  ] = 12'h000;
    rom[256  ] = 12'h000;
    rom[257  ] = 12'h000;
    rom[258  ] = 12'h000;
    rom[259  ] = 12'h000;
    rom[260  ] = 12'h000;
    rom[261  ] = 12'h000;
    rom[262  ] = 12'h000;
    rom[263  ] = 12'h000;
    rom[264  ] = 12'h000;
    rom[265  ] = 12'h000;
    rom[266  ] = 12'h000;
    rom[267  ] = 12'h000;
    rom[268  ] = 12'h000;
    rom[269  ] = 12'h000;
    rom[270  ] = 12'h000;
    rom[271  ] = 12'h000;
    rom[272  ] = 12'h000;
    rom[273  ] = 12'h000;
    rom[274  ] = 12'h000;
    rom[275  ] = 12'h000;
    rom[276  ] = 12'h000;
    rom[277  ] = 12'h000;
    rom[278  ] = 12'h000;
    rom[279  ] = 12'h000;
    rom[280  ] = 12'h000;
    rom[281  ] = 12'h000;
    rom[282  ] = 12'h000;
    rom[283  ] = 12'h000;
    rom[284  ] = 12'h000;
    rom[285  ] = 12'h000;
    rom[286  ] = 12'h000;
    rom[287  ] = 12'h000;
    rom[288  ] = 12'h000;
    rom[289  ] = 12'h000;
    rom[290  ] = 12'h000;
    rom[291  ] = 12'h000;
    rom[292  ] = 12'h000;
    rom[293  ] = 12'h000;
    rom[294  ] = 12'h000;
    rom[295  ] = 12'h000;
    rom[296  ] = 12'h000;
    rom[297  ] = 12'h000;
    rom[298  ] = 12'h000;
    rom[299  ] = 12'h000;
    rom[300  ] = 12'h000;
    rom[301  ] = 12'h000;
    rom[302  ] = 12'h000;
    rom[303  ] = 12'hf90;
    rom[304  ] = 12'hf90;
    rom[305  ] = 12'hf90;
    rom[306  ] = 12'hf90;
    rom[307  ] = 12'hf90;
    rom[308  ] = 12'he90;
    rom[309  ] = 12'he90;
    rom[310  ] = 12'he90;
    rom[311  ] = 12'he90;
    rom[312  ] = 12'he90;
    rom[313  ] = 12'he90;
    rom[314  ] = 12'he90;
    rom[315  ] = 12'he90;
    rom[316  ] = 12'he90;
    rom[317  ] = 12'he90;
    rom[318  ] = 12'he90;
    rom[319  ] = 12'he90;
    rom[320  ] = 12'he90;
    rom[321  ] = 12'he90;
    rom[322  ] = 12'he90;
    rom[323  ] = 12'he90;
    rom[324  ] = 12'he90;
    rom[325  ] = 12'he90;
    rom[326  ] = 12'he90;
    rom[327  ] = 12'he90;
    rom[328  ] = 12'he80;
    rom[329  ] = 12'he80;
    rom[330  ] = 12'he80;
    rom[331  ] = 12'he80;
    rom[332  ] = 12'hd80;
    rom[333  ] = 12'hd80;
    rom[334  ] = 12'hd80;
    rom[335  ] = 12'hd80;
    rom[336  ] = 12'hd80;
    rom[337  ] = 12'hd80;
    rom[338  ] = 12'h000;
    rom[339  ] = 12'h000;
    rom[340  ] = 12'h000;
    rom[341  ] = 12'h000;
    rom[342  ] = 12'h000;
    rom[343  ] = 12'h000;
    rom[344  ] = 12'h000;
    rom[345  ] = 12'h000;
    rom[346  ] = 12'h000;
    rom[347  ] = 12'h000;
    rom[348  ] = 12'h000;
    rom[349  ] = 12'h000;
    rom[350  ] = 12'h000;
    rom[351  ] = 12'h000;
    rom[352  ] = 12'h000;
    rom[353  ] = 12'h000;
    rom[354  ] = 12'h000;
    rom[355  ] = 12'h000;
    rom[356  ] = 12'h000;
    rom[357  ] = 12'h000;
    rom[358  ] = 12'h000;
    rom[359  ] = 12'h000;
    rom[360  ] = 12'h000;
    rom[361  ] = 12'h000;
    rom[362  ] = 12'h000;
    rom[363  ] = 12'h000;
    rom[364  ] = 12'h000;
    rom[365  ] = 12'h000;
    rom[366  ] = 12'h000;
    rom[367  ] = 12'h000;
    rom[368  ] = 12'h000;
    rom[369  ] = 12'h000;
    rom[370  ] = 12'h000;
    rom[371  ] = 12'h000;
    rom[372  ] = 12'h000;
    rom[373  ] = 12'h000;
    rom[374  ] = 12'h000;
    rom[375  ] = 12'h000;
    rom[376  ] = 12'h000;
    rom[377  ] = 12'h000;
    rom[378  ] = 12'h000;
    rom[379  ] = 12'h000;
    rom[380  ] = 12'h000;
    rom[381  ] = 12'h000;
    rom[382  ] = 12'h000;
    rom[383  ] = 12'h000;
    rom[384  ] = 12'h000;
    rom[385  ] = 12'h000;
    rom[386  ] = 12'h000;
    rom[387  ] = 12'h000;
    rom[388  ] = 12'h000;
    rom[389  ] = 12'h000;
    rom[390  ] = 12'h000;
    rom[391  ] = 12'h000;
    rom[392  ] = 12'h000;
    rom[393  ] = 12'h000;
    rom[394  ] = 12'h000;
    rom[395  ] = 12'h000;
    rom[396  ] = 12'h000;
    rom[397  ] = 12'h000;
    rom[398  ] = 12'h000;
    rom[399  ] = 12'h000;
    rom[400  ] = 12'h000;
    rom[401  ] = 12'h000;
    rom[402  ] = 12'h000;
    rom[403  ] = 12'h000;
    rom[404  ] = 12'h000;
    rom[405  ] = 12'h000;
    rom[406  ] = 12'h000;
    rom[407  ] = 12'h000;
    rom[408  ] = 12'h000;
    rom[409  ] = 12'h000;
    rom[410  ] = 12'h000;
    rom[411  ] = 12'h000;
    rom[412  ] = 12'h000;
    rom[413  ] = 12'h000;
    rom[414  ] = 12'h000;
    rom[415  ] = 12'h000;
    rom[416  ] = 12'h000;
    rom[417  ] = 12'h000;
    rom[418  ] = 12'h000;
    rom[419  ] = 12'h000;
    rom[420  ] = 12'h000;
    rom[421  ] = 12'h000;
    rom[422  ] = 12'h000;
    rom[423  ] = 12'h000;
    rom[424  ] = 12'h000;
    rom[425  ] = 12'h000;
    rom[426  ] = 12'h000;
    rom[427  ] = 12'hf90;
    rom[428  ] = 12'hf90;
    rom[429  ] = 12'hf90;
    rom[430  ] = 12'hf90;
    rom[431  ] = 12'hf90;
    rom[432  ] = 12'hf90;
    rom[433  ] = 12'hf90;
    rom[434  ] = 12'hf90;
    rom[435  ] = 12'hf90;
    rom[436  ] = 12'hf90;
    rom[437  ] = 12'he90;
    rom[438  ] = 12'he90;
    rom[439  ] = 12'he90;
    rom[440  ] = 12'he90;
    rom[441  ] = 12'he90;
    rom[442  ] = 12'he90;
    rom[443  ] = 12'he90;
    rom[444  ] = 12'he90;
    rom[445  ] = 12'he90;
    rom[446  ] = 12'he90;
    rom[447  ] = 12'he90;
    rom[448  ] = 12'he90;
    rom[449  ] = 12'he90;
    rom[450  ] = 12'he90;
    rom[451  ] = 12'he90;
    rom[452  ] = 12'he90;
    rom[453  ] = 12'he90;
    rom[454  ] = 12'he90;
    rom[455  ] = 12'he90;
    rom[456  ] = 12'he80;
    rom[457  ] = 12'he80;
    rom[458  ] = 12'he80;
    rom[459  ] = 12'he80;
    rom[460  ] = 12'hd80;
    rom[461  ] = 12'hd80;
    rom[462  ] = 12'hd80;
    rom[463  ] = 12'hd80;
    rom[464  ] = 12'hd80;
    rom[465  ] = 12'hd80;
    rom[466  ] = 12'hd80;
    rom[467  ] = 12'hd80;
    rom[468  ] = 12'hd80;
    rom[469  ] = 12'h000;
    rom[470  ] = 12'h000;
    rom[471  ] = 12'h000;
    rom[472  ] = 12'h000;
    rom[473  ] = 12'h000;
    rom[474  ] = 12'h000;
    rom[475  ] = 12'h000;
    rom[476  ] = 12'h000;
    rom[477  ] = 12'h000;
    rom[478  ] = 12'h000;
    rom[479  ] = 12'h000;
    rom[480  ] = 12'h000;
    rom[481  ] = 12'h000;
    rom[482  ] = 12'h000;
    rom[483  ] = 12'h000;
    rom[484  ] = 12'h000;
    rom[485  ] = 12'h000;
    rom[486  ] = 12'h000;
    rom[487  ] = 12'h000;
    rom[488  ] = 12'h000;
    rom[489  ] = 12'h000;
    rom[490  ] = 12'h000;
    rom[491  ] = 12'h000;
    rom[492  ] = 12'h000;
    rom[493  ] = 12'h000;
    rom[494  ] = 12'h000;
    rom[495  ] = 12'h000;
    rom[496  ] = 12'h000;
    rom[497  ] = 12'h000;
    rom[498  ] = 12'h000;
    rom[499  ] = 12'h000;
    rom[500  ] = 12'h000;
    rom[501  ] = 12'h000;
    rom[502  ] = 12'h000;
    rom[503  ] = 12'h000;
    rom[504  ] = 12'h000;
    rom[505  ] = 12'h000;
    rom[506  ] = 12'h000;
    rom[507  ] = 12'h000;
    rom[508  ] = 12'h000;
    rom[509  ] = 12'h000;
    rom[510  ] = 12'h000;
    rom[511  ] = 12'h000;
    rom[512  ] = 12'h000;
    rom[513  ] = 12'h000;
    rom[514  ] = 12'h000;
    rom[515  ] = 12'h000;
    rom[516  ] = 12'h000;
    rom[517  ] = 12'h000;
    rom[518  ] = 12'h000;
    rom[519  ] = 12'h000;
    rom[520  ] = 12'h000;
    rom[521  ] = 12'h000;
    rom[522  ] = 12'h000;
    rom[523  ] = 12'h000;
    rom[524  ] = 12'h000;
    rom[525  ] = 12'h000;
    rom[526  ] = 12'h000;
    rom[527  ] = 12'h000;
    rom[528  ] = 12'h000;
    rom[529  ] = 12'h000;
    rom[530  ] = 12'h000;
    rom[531  ] = 12'h000;
    rom[532  ] = 12'h000;
    rom[533  ] = 12'h000;
    rom[534  ] = 12'h000;
    rom[535  ] = 12'h000;
    rom[536  ] = 12'h000;
    rom[537  ] = 12'h000;
    rom[538  ] = 12'h000;
    rom[539  ] = 12'h000;
    rom[540  ] = 12'h000;
    rom[541  ] = 12'h000;
    rom[542  ] = 12'h000;
    rom[543  ] = 12'h000;
    rom[544  ] = 12'h000;
    rom[545  ] = 12'h000;
    rom[546  ] = 12'h000;
    rom[547  ] = 12'h000;
    rom[548  ] = 12'h000;
    rom[549  ] = 12'h000;
    rom[550  ] = 12'h000;
    rom[551  ] = 12'h000;
    rom[552  ] = 12'h000;
    rom[553  ] = 12'hf90;
    rom[554  ] = 12'hf90;
    rom[555  ] = 12'hf90;
    rom[556  ] = 12'hf90;
    rom[557  ] = 12'hf90;
    rom[558  ] = 12'hf90;
    rom[559  ] = 12'hf90;
    rom[560  ] = 12'hf90;
    rom[561  ] = 12'hf90;
    rom[562  ] = 12'hf90;
    rom[563  ] = 12'hf90;
    rom[564  ] = 12'hf90;
    rom[565  ] = 12'he90;
    rom[566  ] = 12'he90;
    rom[567  ] = 12'he90;
    rom[568  ] = 12'he90;
    rom[569  ] = 12'he90;
    rom[570  ] = 12'he90;
    rom[571  ] = 12'he90;
    rom[572  ] = 12'he90;
    rom[573  ] = 12'he90;
    rom[574  ] = 12'he90;
    rom[575  ] = 12'he90;
    rom[576  ] = 12'he90;
    rom[577  ] = 12'he90;
    rom[578  ] = 12'he90;
    rom[579  ] = 12'he90;
    rom[580  ] = 12'he90;
    rom[581  ] = 12'he90;
    rom[582  ] = 12'he90;
    rom[583  ] = 12'he80;
    rom[584  ] = 12'he80;
    rom[585  ] = 12'he80;
    rom[586  ] = 12'he80;
    rom[587  ] = 12'he80;
    rom[588  ] = 12'hd80;
    rom[589  ] = 12'hd80;
    rom[590  ] = 12'hd80;
    rom[591  ] = 12'hd80;
    rom[592  ] = 12'hd80;
    rom[593  ] = 12'hd80;
    rom[594  ] = 12'hd80;
    rom[595  ] = 12'hd80;
    rom[596  ] = 12'hd80;
    rom[597  ] = 12'hd80;
    rom[598  ] = 12'hd80;
    rom[599  ] = 12'h000;
    rom[600  ] = 12'h000;
    rom[601  ] = 12'h000;
    rom[602  ] = 12'h000;
    rom[603  ] = 12'h000;
    rom[604  ] = 12'h000;
    rom[605  ] = 12'h000;
    rom[606  ] = 12'h000;
    rom[607  ] = 12'h000;
    rom[608  ] = 12'h000;
    rom[609  ] = 12'h000;
    rom[610  ] = 12'h000;
    rom[611  ] = 12'h000;
    rom[612  ] = 12'h000;
    rom[613  ] = 12'h000;
    rom[614  ] = 12'h000;
    rom[615  ] = 12'h000;
    rom[616  ] = 12'h000;
    rom[617  ] = 12'h000;
    rom[618  ] = 12'h000;
    rom[619  ] = 12'h000;
    rom[620  ] = 12'h000;
    rom[621  ] = 12'h000;
    rom[622  ] = 12'h000;
    rom[623  ] = 12'h000;
    rom[624  ] = 12'h000;
    rom[625  ] = 12'h000;
    rom[626  ] = 12'h000;
    rom[627  ] = 12'h000;
    rom[628  ] = 12'h000;
    rom[629  ] = 12'h000;
    rom[630  ] = 12'h000;
    rom[631  ] = 12'h000;
    rom[632  ] = 12'h000;
    rom[633  ] = 12'h000;
    rom[634  ] = 12'h000;
    rom[635  ] = 12'h000;
    rom[636  ] = 12'h000;
    rom[637  ] = 12'h000;
    rom[638  ] = 12'h000;
    rom[639  ] = 12'h000;
    rom[640  ] = 12'h000;
    rom[641  ] = 12'h000;
    rom[642  ] = 12'h000;
    rom[643  ] = 12'h000;
    rom[644  ] = 12'h000;
    rom[645  ] = 12'h000;
    rom[646  ] = 12'h000;
    rom[647  ] = 12'h000;
    rom[648  ] = 12'h000;
    rom[649  ] = 12'h000;
    rom[650  ] = 12'h000;
    rom[651  ] = 12'h000;
    rom[652  ] = 12'h000;
    rom[653  ] = 12'h000;
    rom[654  ] = 12'h000;
    rom[655  ] = 12'h000;
    rom[656  ] = 12'h000;
    rom[657  ] = 12'h000;
    rom[658  ] = 12'h000;
    rom[659  ] = 12'h000;
    rom[660  ] = 12'h000;
    rom[661  ] = 12'h000;
    rom[662  ] = 12'h000;
    rom[663  ] = 12'h000;
    rom[664  ] = 12'h000;
    rom[665  ] = 12'h000;
    rom[666  ] = 12'h000;
    rom[667  ] = 12'h000;
    rom[668  ] = 12'h000;
    rom[669  ] = 12'h000;
    rom[670  ] = 12'h000;
    rom[671  ] = 12'h000;
    rom[672  ] = 12'h000;
    rom[673  ] = 12'h000;
    rom[674  ] = 12'h000;
    rom[675  ] = 12'h000;
    rom[676  ] = 12'h000;
    rom[677  ] = 12'h000;
    rom[678  ] = 12'hf90;
    rom[679  ] = 12'hf90;
    rom[680  ] = 12'hf90;
    rom[681  ] = 12'hf90;
    rom[682  ] = 12'hf90;
    rom[683  ] = 12'hf90;
    rom[684  ] = 12'hf90;
    rom[685  ] = 12'hf90;
    rom[686  ] = 12'hf90;
    rom[687  ] = 12'hf90;
    rom[688  ] = 12'hf90;
    rom[689  ] = 12'hf90;
    rom[690  ] = 12'hf90;
    rom[691  ] = 12'hf90;
    rom[692  ] = 12'hf90;
    rom[693  ] = 12'he90;
    rom[694  ] = 12'he90;
    rom[695  ] = 12'he90;
    rom[696  ] = 12'he90;
    rom[697  ] = 12'he90;
    rom[698  ] = 12'he90;
    rom[699  ] = 12'he90;
    rom[700  ] = 12'he90;
    rom[701  ] = 12'he90;
    rom[702  ] = 12'he90;
    rom[703  ] = 12'he90;
    rom[704  ] = 12'he90;
    rom[705  ] = 12'he90;
    rom[706  ] = 12'he90;
    rom[707  ] = 12'he90;
    rom[708  ] = 12'he90;
    rom[709  ] = 12'he90;
    rom[710  ] = 12'he90;
    rom[711  ] = 12'he80;
    rom[712  ] = 12'he80;
    rom[713  ] = 12'he80;
    rom[714  ] = 12'he80;
    rom[715  ] = 12'hd80;
    rom[716  ] = 12'hd80;
    rom[717  ] = 12'hd80;
    rom[718  ] = 12'hd80;
    rom[719  ] = 12'hd80;
    rom[720  ] = 12'hd80;
    rom[721  ] = 12'hd80;
    rom[722  ] = 12'hd80;
    rom[723  ] = 12'hd80;
    rom[724  ] = 12'hd80;
    rom[725  ] = 12'hd80;
    rom[726  ] = 12'hd80;
    rom[727  ] = 12'hd80;
    rom[728  ] = 12'hd80;
    rom[729  ] = 12'hd80;
    rom[730  ] = 12'h000;
    rom[731  ] = 12'h000;
    rom[732  ] = 12'h000;
    rom[733  ] = 12'h000;
    rom[734  ] = 12'h000;
    rom[735  ] = 12'h000;
    rom[736  ] = 12'h000;
    rom[737  ] = 12'h000;
    rom[738  ] = 12'h000;
    rom[739  ] = 12'h000;
    rom[740  ] = 12'h000;
    rom[741  ] = 12'h000;
    rom[742  ] = 12'h000;
    rom[743  ] = 12'h000;
    rom[744  ] = 12'h000;
    rom[745  ] = 12'h000;
    rom[746  ] = 12'h000;
    rom[747  ] = 12'h000;
    rom[748  ] = 12'h000;
    rom[749  ] = 12'h000;
    rom[750  ] = 12'h000;
    rom[751  ] = 12'h000;
    rom[752  ] = 12'h000;
    rom[753  ] = 12'h000;
    rom[754  ] = 12'h000;
    rom[755  ] = 12'h000;
    rom[756  ] = 12'h000;
    rom[757  ] = 12'h000;
    rom[758  ] = 12'h000;
    rom[759  ] = 12'h000;
    rom[760  ] = 12'h000;
    rom[761  ] = 12'h000;
    rom[762  ] = 12'h000;
    rom[763  ] = 12'h000;
    rom[764  ] = 12'h000;
    rom[765  ] = 12'h000;
    rom[766  ] = 12'h000;
    rom[767  ] = 12'h000;
    rom[768  ] = 12'h000;
    rom[769  ] = 12'h000;
    rom[770  ] = 12'h000;
    rom[771  ] = 12'h000;
    rom[772  ] = 12'h000;
    rom[773  ] = 12'h000;
    rom[774  ] = 12'h000;
    rom[775  ] = 12'h000;
    rom[776  ] = 12'h000;
    rom[777  ] = 12'h000;
    rom[778  ] = 12'h000;
    rom[779  ] = 12'h000;
    rom[780  ] = 12'h000;
    rom[781  ] = 12'h000;
    rom[782  ] = 12'h000;
    rom[783  ] = 12'h000;
    rom[784  ] = 12'h000;
    rom[785  ] = 12'h000;
    rom[786  ] = 12'h000;
    rom[787  ] = 12'h000;
    rom[788  ] = 12'h000;
    rom[789  ] = 12'h000;
    rom[790  ] = 12'h000;
    rom[791  ] = 12'h000;
    rom[792  ] = 12'h000;
    rom[793  ] = 12'h000;
    rom[794  ] = 12'h000;
    rom[795  ] = 12'h000;
    rom[796  ] = 12'h000;
    rom[797  ] = 12'h000;
    rom[798  ] = 12'h000;
    rom[799  ] = 12'h000;
    rom[800  ] = 12'h000;
    rom[801  ] = 12'h000;
    rom[802  ] = 12'h000;
    rom[803  ] = 12'h000;
    rom[804  ] = 12'hf90;
    rom[805  ] = 12'hf90;
    rom[806  ] = 12'hf90;
    rom[807  ] = 12'hf90;
    rom[808  ] = 12'hf90;
    rom[809  ] = 12'hf90;
    rom[810  ] = 12'hf90;
    rom[811  ] = 12'hf90;
    rom[812  ] = 12'hf90;
    rom[813  ] = 12'hf90;
    rom[814  ] = 12'hf90;
    rom[815  ] = 12'hf90;
    rom[816  ] = 12'hf90;
    rom[817  ] = 12'hf90;
    rom[818  ] = 12'hf90;
    rom[819  ] = 12'hf90;
    rom[820  ] = 12'hf90;
    rom[821  ] = 12'hf90;
    rom[822  ] = 12'he90;
    rom[823  ] = 12'he90;
    rom[824  ] = 12'he90;
    rom[825  ] = 12'he90;
    rom[826  ] = 12'he90;
    rom[827  ] = 12'he90;
    rom[828  ] = 12'he90;
    rom[829  ] = 12'he90;
    rom[830  ] = 12'he90;
    rom[831  ] = 12'he90;
    rom[832  ] = 12'he90;
    rom[833  ] = 12'he90;
    rom[834  ] = 12'he90;
    rom[835  ] = 12'he90;
    rom[836  ] = 12'he90;
    rom[837  ] = 12'he90;
    rom[838  ] = 12'he90;
    rom[839  ] = 12'he80;
    rom[840  ] = 12'he80;
    rom[841  ] = 12'he80;
    rom[842  ] = 12'he80;
    rom[843  ] = 12'hd80;
    rom[844  ] = 12'hd80;
    rom[845  ] = 12'hd80;
    rom[846  ] = 12'hd80;
    rom[847  ] = 12'hd80;
    rom[848  ] = 12'hd80;
    rom[849  ] = 12'hd80;
    rom[850  ] = 12'hd80;
    rom[851  ] = 12'hd80;
    rom[852  ] = 12'hd80;
    rom[853  ] = 12'hd80;
    rom[854  ] = 12'hd80;
    rom[855  ] = 12'hd80;
    rom[856  ] = 12'hd80;
    rom[857  ] = 12'hd80;
    rom[858  ] = 12'hc80;
    rom[859  ] = 12'hc80;
    rom[860  ] = 12'h000;
    rom[861  ] = 12'h000;
    rom[862  ] = 12'h000;
    rom[863  ] = 12'h000;
    rom[864  ] = 12'h000;
    rom[865  ] = 12'h000;
    rom[866  ] = 12'h000;
    rom[867  ] = 12'h000;
    rom[868  ] = 12'h000;
    rom[869  ] = 12'h000;
    rom[870  ] = 12'h000;
    rom[871  ] = 12'h000;
    rom[872  ] = 12'h000;
    rom[873  ] = 12'h000;
    rom[874  ] = 12'h000;
    rom[875  ] = 12'h000;
    rom[876  ] = 12'h000;
    rom[877  ] = 12'h000;
    rom[878  ] = 12'h000;
    rom[879  ] = 12'h000;
    rom[880  ] = 12'h000;
    rom[881  ] = 12'h000;
    rom[882  ] = 12'h000;
    rom[883  ] = 12'h000;
    rom[884  ] = 12'h000;
    rom[885  ] = 12'h000;
    rom[886  ] = 12'h000;
    rom[887  ] = 12'h000;
    rom[888  ] = 12'h000;
    rom[889  ] = 12'h000;
    rom[890  ] = 12'h000;
    rom[891  ] = 12'h000;
    rom[892  ] = 12'h000;
    rom[893  ] = 12'h000;
    rom[894  ] = 12'h000;
    rom[895  ] = 12'h000;
    rom[896  ] = 12'h000;
    rom[897  ] = 12'h000;
    rom[898  ] = 12'h000;
    rom[899  ] = 12'h000;
    rom[900  ] = 12'h000;
    rom[901  ] = 12'h000;
    rom[902  ] = 12'h000;
    rom[903  ] = 12'h000;
    rom[904  ] = 12'h000;
    rom[905  ] = 12'h000;
    rom[906  ] = 12'h000;
    rom[907  ] = 12'h000;
    rom[908  ] = 12'h000;
    rom[909  ] = 12'h000;
    rom[910  ] = 12'h000;
    rom[911  ] = 12'h000;
    rom[912  ] = 12'h000;
    rom[913  ] = 12'h000;
    rom[914  ] = 12'h000;
    rom[915  ] = 12'h000;
    rom[916  ] = 12'h000;
    rom[917  ] = 12'h000;
    rom[918  ] = 12'h000;
    rom[919  ] = 12'h000;
    rom[920  ] = 12'h000;
    rom[921  ] = 12'h000;
    rom[922  ] = 12'h000;
    rom[923  ] = 12'h000;
    rom[924  ] = 12'h000;
    rom[925  ] = 12'h000;
    rom[926  ] = 12'h000;
    rom[927  ] = 12'h000;
    rom[928  ] = 12'h000;
    rom[929  ] = 12'h000;
    rom[930  ] = 12'he90;
    rom[931  ] = 12'hf90;
    rom[932  ] = 12'hf90;
    rom[933  ] = 12'hf90;
    rom[934  ] = 12'hf90;
    rom[935  ] = 12'hf90;
    rom[936  ] = 12'hf90;
    rom[937  ] = 12'hf90;
    rom[938  ] = 12'hf90;
    rom[939  ] = 12'hf90;
    rom[940  ] = 12'hf90;
    rom[941  ] = 12'hf90;
    rom[942  ] = 12'hf90;
    rom[943  ] = 12'hf90;
    rom[944  ] = 12'hf90;
    rom[945  ] = 12'hf90;
    rom[946  ] = 12'hf90;
    rom[947  ] = 12'hf90;
    rom[948  ] = 12'hf90;
    rom[949  ] = 12'hf90;
    rom[950  ] = 12'he90;
    rom[951  ] = 12'he90;
    rom[952  ] = 12'he90;
    rom[953  ] = 12'he90;
    rom[954  ] = 12'he90;
    rom[955  ] = 12'he90;
    rom[956  ] = 12'he90;
    rom[957  ] = 12'he90;
    rom[958  ] = 12'he90;
    rom[959  ] = 12'he90;
    rom[960  ] = 12'he90;
    rom[961  ] = 12'he90;
    rom[962  ] = 12'he90;
    rom[963  ] = 12'he90;
    rom[964  ] = 12'he90;
    rom[965  ] = 12'he90;
    rom[966  ] = 12'he80;
    rom[967  ] = 12'he80;
    rom[968  ] = 12'he80;
    rom[969  ] = 12'he80;
    rom[970  ] = 12'he80;
    rom[971  ] = 12'hd80;
    rom[972  ] = 12'hd80;
    rom[973  ] = 12'hd80;
    rom[974  ] = 12'hd80;
    rom[975  ] = 12'hd80;
    rom[976  ] = 12'hd80;
    rom[977  ] = 12'hd80;
    rom[978  ] = 12'hd80;
    rom[979  ] = 12'hd80;
    rom[980  ] = 12'hd80;
    rom[981  ] = 12'hd80;
    rom[982  ] = 12'hd80;
    rom[983  ] = 12'hd80;
    rom[984  ] = 12'hd80;
    rom[985  ] = 12'hd80;
    rom[986  ] = 12'hc80;
    rom[987  ] = 12'hc80;
    rom[988  ] = 12'hc80;
    rom[989  ] = 12'hc80;
    rom[990  ] = 12'h000;
    rom[991  ] = 12'h000;
    rom[992  ] = 12'h000;
    rom[993  ] = 12'h000;
    rom[994  ] = 12'h000;
    rom[995  ] = 12'h000;
    rom[996  ] = 12'h000;
    rom[997  ] = 12'h000;
    rom[998  ] = 12'h000;
    rom[999  ] = 12'h000;
    rom[1000 ] = 12'h000;
    rom[1001 ] = 12'h000;
    rom[1002 ] = 12'h000;
    rom[1003 ] = 12'h000;
    rom[1004 ] = 12'h000;
    rom[1005 ] = 12'h000;
    rom[1006 ] = 12'h000;
    rom[1007 ] = 12'h000;
    rom[1008 ] = 12'h000;
    rom[1009 ] = 12'h000;
    rom[1010 ] = 12'h000;
    rom[1011 ] = 12'h000;
    rom[1012 ] = 12'h000;
    rom[1013 ] = 12'h000;
    rom[1014 ] = 12'h000;
    rom[1015 ] = 12'h000;
    rom[1016 ] = 12'h000;
    rom[1017 ] = 12'h000;
    rom[1018 ] = 12'h000;
    rom[1019 ] = 12'h000;
    rom[1020 ] = 12'h000;
    rom[1021 ] = 12'h000;
    rom[1022 ] = 12'h000;
    rom[1023 ] = 12'h000;
    rom[1024 ] = 12'h000;
    rom[1025 ] = 12'h000;
    rom[1026 ] = 12'h000;
    rom[1027 ] = 12'h000;
    rom[1028 ] = 12'h000;
    rom[1029 ] = 12'h000;
    rom[1030 ] = 12'h000;
    rom[1031 ] = 12'h000;
    rom[1032 ] = 12'h000;
    rom[1033 ] = 12'h000;
    rom[1034 ] = 12'h000;
    rom[1035 ] = 12'h000;
    rom[1036 ] = 12'h000;
    rom[1037 ] = 12'h000;
    rom[1038 ] = 12'h000;
    rom[1039 ] = 12'h000;
    rom[1040 ] = 12'h000;
    rom[1041 ] = 12'h000;
    rom[1042 ] = 12'h000;
    rom[1043 ] = 12'h000;
    rom[1044 ] = 12'h000;
    rom[1045 ] = 12'h000;
    rom[1046 ] = 12'h000;
    rom[1047 ] = 12'h000;
    rom[1048 ] = 12'h000;
    rom[1049 ] = 12'h000;
    rom[1050 ] = 12'h000;
    rom[1051 ] = 12'h000;
    rom[1052 ] = 12'h000;
    rom[1053 ] = 12'h000;
    rom[1054 ] = 12'h000;
    rom[1055 ] = 12'h000;
    rom[1056 ] = 12'hea0;
    rom[1057 ] = 12'hea0;
    rom[1058 ] = 12'he90;
    rom[1059 ] = 12'hf90;
    rom[1060 ] = 12'hf90;
    rom[1061 ] = 12'hf90;
    rom[1062 ] = 12'hf90;
    rom[1063 ] = 12'hf90;
    rom[1064 ] = 12'hf90;
    rom[1065 ] = 12'hf90;
    rom[1066 ] = 12'hf90;
    rom[1067 ] = 12'hf90;
    rom[1068 ] = 12'hf90;
    rom[1069 ] = 12'hf90;
    rom[1070 ] = 12'hf90;
    rom[1071 ] = 12'hf90;
    rom[1072 ] = 12'hf90;
    rom[1073 ] = 12'hf90;
    rom[1074 ] = 12'hf90;
    rom[1075 ] = 12'hf90;
    rom[1076 ] = 12'hf90;
    rom[1077 ] = 12'hf90;
    rom[1078 ] = 12'hf90;
    rom[1079 ] = 12'he90;
    rom[1080 ] = 12'he90;
    rom[1081 ] = 12'he90;
    rom[1082 ] = 12'he90;
    rom[1083 ] = 12'he90;
    rom[1084 ] = 12'he90;
    rom[1085 ] = 12'he90;
    rom[1086 ] = 12'he90;
    rom[1087 ] = 12'he90;
    rom[1088 ] = 12'he90;
    rom[1089 ] = 12'he90;
    rom[1090 ] = 12'he90;
    rom[1091 ] = 12'he90;
    rom[1092 ] = 12'he90;
    rom[1093 ] = 12'he90;
    rom[1094 ] = 12'he80;
    rom[1095 ] = 12'he80;
    rom[1096 ] = 12'he80;
    rom[1097 ] = 12'he80;
    rom[1098 ] = 12'hd80;
    rom[1099 ] = 12'hd80;
    rom[1100 ] = 12'hd80;
    rom[1101 ] = 12'hd80;
    rom[1102 ] = 12'hd80;
    rom[1103 ] = 12'hd80;
    rom[1104 ] = 12'hd80;
    rom[1105 ] = 12'hd80;
    rom[1106 ] = 12'hd80;
    rom[1107 ] = 12'hd80;
    rom[1108 ] = 12'hd80;
    rom[1109 ] = 12'hd80;
    rom[1110 ] = 12'hd80;
    rom[1111 ] = 12'hd80;
    rom[1112 ] = 12'hd80;
    rom[1113 ] = 12'hd80;
    rom[1114 ] = 12'hc80;
    rom[1115 ] = 12'hc80;
    rom[1116 ] = 12'hc80;
    rom[1117 ] = 12'hc80;
    rom[1118 ] = 12'hc80;
    rom[1119 ] = 12'hc80;
    rom[1120 ] = 12'h000;
    rom[1121 ] = 12'h000;
    rom[1122 ] = 12'h000;
    rom[1123 ] = 12'h000;
    rom[1124 ] = 12'h000;
    rom[1125 ] = 12'h000;
    rom[1126 ] = 12'h000;
    rom[1127 ] = 12'h000;
    rom[1128 ] = 12'h000;
    rom[1129 ] = 12'h000;
    rom[1130 ] = 12'h000;
    rom[1131 ] = 12'h000;
    rom[1132 ] = 12'h000;
    rom[1133 ] = 12'h000;
    rom[1134 ] = 12'h000;
    rom[1135 ] = 12'h000;
    rom[1136 ] = 12'h000;
    rom[1137 ] = 12'h000;
    rom[1138 ] = 12'h000;
    rom[1139 ] = 12'h000;
    rom[1140 ] = 12'h000;
    rom[1141 ] = 12'h000;
    rom[1142 ] = 12'h000;
    rom[1143 ] = 12'h000;
    rom[1144 ] = 12'h000;
    rom[1145 ] = 12'h000;
    rom[1146 ] = 12'h000;
    rom[1147 ] = 12'h000;
    rom[1148 ] = 12'h000;
    rom[1149 ] = 12'h000;
    rom[1150 ] = 12'h000;
    rom[1151 ] = 12'h000;
    rom[1152 ] = 12'h000;
    rom[1153 ] = 12'h000;
    rom[1154 ] = 12'h000;
    rom[1155 ] = 12'h000;
    rom[1156 ] = 12'h000;
    rom[1157 ] = 12'h000;
    rom[1158 ] = 12'h000;
    rom[1159 ] = 12'h000;
    rom[1160 ] = 12'h000;
    rom[1161 ] = 12'h000;
    rom[1162 ] = 12'h000;
    rom[1163 ] = 12'h000;
    rom[1164 ] = 12'h000;
    rom[1165 ] = 12'h000;
    rom[1166 ] = 12'h000;
    rom[1167 ] = 12'h000;
    rom[1168 ] = 12'h000;
    rom[1169 ] = 12'h000;
    rom[1170 ] = 12'h000;
    rom[1171 ] = 12'h000;
    rom[1172 ] = 12'h000;
    rom[1173 ] = 12'h000;
    rom[1174 ] = 12'h000;
    rom[1175 ] = 12'h000;
    rom[1176 ] = 12'h000;
    rom[1177 ] = 12'h000;
    rom[1178 ] = 12'h000;
    rom[1179 ] = 12'h000;
    rom[1180 ] = 12'h000;
    rom[1181 ] = 12'h000;
    rom[1182 ] = 12'h000;
    rom[1183 ] = 12'hea0;
    rom[1184 ] = 12'hea0;
    rom[1185 ] = 12'hea0;
    rom[1186 ] = 12'hea0;
    rom[1187 ] = 12'he90;
    rom[1188 ] = 12'hf90;
    rom[1189 ] = 12'hf90;
    rom[1190 ] = 12'hf90;
    rom[1191 ] = 12'hf90;
    rom[1192 ] = 12'hf90;
    rom[1193 ] = 12'hf90;
    rom[1194 ] = 12'hf90;
    rom[1195 ] = 12'hf90;
    rom[1196 ] = 12'hf90;
    rom[1197 ] = 12'hf90;
    rom[1198 ] = 12'hf90;
    rom[1199 ] = 12'hf90;
    rom[1200 ] = 12'hf90;
    rom[1201 ] = 12'hf90;
    rom[1202 ] = 12'hf90;
    rom[1203 ] = 12'hf90;
    rom[1204 ] = 12'hf90;
    rom[1205 ] = 12'hf90;
    rom[1206 ] = 12'hf90;
    rom[1207 ] = 12'he90;
    rom[1208 ] = 12'he90;
    rom[1209 ] = 12'he90;
    rom[1210 ] = 12'he90;
    rom[1211 ] = 12'he90;
    rom[1212 ] = 12'he90;
    rom[1213 ] = 12'he90;
    rom[1214 ] = 12'he90;
    rom[1215 ] = 12'he90;
    rom[1216 ] = 12'he90;
    rom[1217 ] = 12'he90;
    rom[1218 ] = 12'he90;
    rom[1219 ] = 12'he90;
    rom[1220 ] = 12'he90;
    rom[1221 ] = 12'he90;
    rom[1222 ] = 12'he80;
    rom[1223 ] = 12'he80;
    rom[1224 ] = 12'he80;
    rom[1225 ] = 12'he80;
    rom[1226 ] = 12'hd80;
    rom[1227 ] = 12'hd80;
    rom[1228 ] = 12'hd80;
    rom[1229 ] = 12'hd80;
    rom[1230 ] = 12'hd80;
    rom[1231 ] = 12'hd80;
    rom[1232 ] = 12'hd80;
    rom[1233 ] = 12'hd80;
    rom[1234 ] = 12'hd80;
    rom[1235 ] = 12'hd80;
    rom[1236 ] = 12'hd80;
    rom[1237 ] = 12'hd80;
    rom[1238 ] = 12'hd80;
    rom[1239 ] = 12'hd80;
    rom[1240 ] = 12'hd80;
    rom[1241 ] = 12'hc80;
    rom[1242 ] = 12'hc80;
    rom[1243 ] = 12'hc80;
    rom[1244 ] = 12'hc80;
    rom[1245 ] = 12'hc80;
    rom[1246 ] = 12'hc80;
    rom[1247 ] = 12'hc80;
    rom[1248 ] = 12'hc80;
    rom[1249 ] = 12'h000;
    rom[1250 ] = 12'h000;
    rom[1251 ] = 12'h000;
    rom[1252 ] = 12'h000;
    rom[1253 ] = 12'h000;
    rom[1254 ] = 12'h000;
    rom[1255 ] = 12'h000;
    rom[1256 ] = 12'h000;
    rom[1257 ] = 12'h000;
    rom[1258 ] = 12'h000;
    rom[1259 ] = 12'h000;
    rom[1260 ] = 12'h000;
    rom[1261 ] = 12'h000;
    rom[1262 ] = 12'h000;
    rom[1263 ] = 12'h000;
    rom[1264 ] = 12'h000;
    rom[1265 ] = 12'h000;
    rom[1266 ] = 12'h000;
    rom[1267 ] = 12'h000;
    rom[1268 ] = 12'h000;
    rom[1269 ] = 12'h000;
    rom[1270 ] = 12'h000;
    rom[1271 ] = 12'h000;
    rom[1272 ] = 12'h000;
    rom[1273 ] = 12'h000;
    rom[1274 ] = 12'h000;
    rom[1275 ] = 12'h000;
    rom[1276 ] = 12'h000;
    rom[1277 ] = 12'h000;
    rom[1278 ] = 12'h000;
    rom[1279 ] = 12'h000;
    rom[1280 ] = 12'h000;
    rom[1281 ] = 12'h000;
    rom[1282 ] = 12'h000;
    rom[1283 ] = 12'h000;
    rom[1284 ] = 12'h000;
    rom[1285 ] = 12'h000;
    rom[1286 ] = 12'h000;
    rom[1287 ] = 12'h000;
    rom[1288 ] = 12'h000;
    rom[1289 ] = 12'h000;
    rom[1290 ] = 12'h000;
    rom[1291 ] = 12'h000;
    rom[1292 ] = 12'h000;
    rom[1293 ] = 12'h000;
    rom[1294 ] = 12'h000;
    rom[1295 ] = 12'h000;
    rom[1296 ] = 12'h000;
    rom[1297 ] = 12'h000;
    rom[1298 ] = 12'h000;
    rom[1299 ] = 12'h000;
    rom[1300 ] = 12'h000;
    rom[1301 ] = 12'h000;
    rom[1302 ] = 12'h000;
    rom[1303 ] = 12'h000;
    rom[1304 ] = 12'h000;
    rom[1305 ] = 12'h000;
    rom[1306 ] = 12'h000;
    rom[1307 ] = 12'h000;
    rom[1308 ] = 12'h000;
    rom[1309 ] = 12'hea0;
    rom[1310 ] = 12'hea0;
    rom[1311 ] = 12'hea0;
    rom[1312 ] = 12'hea0;
    rom[1313 ] = 12'hea0;
    rom[1314 ] = 12'hea0;
    rom[1315 ] = 12'he90;
    rom[1316 ] = 12'hf90;
    rom[1317 ] = 12'hf90;
    rom[1318 ] = 12'hf90;
    rom[1319 ] = 12'hf90;
    rom[1320 ] = 12'hf90;
    rom[1321 ] = 12'hf90;
    rom[1322 ] = 12'hf90;
    rom[1323 ] = 12'hf90;
    rom[1324 ] = 12'hf90;
    rom[1325 ] = 12'hf90;
    rom[1326 ] = 12'hf90;
    rom[1327 ] = 12'hf90;
    rom[1328 ] = 12'hf90;
    rom[1329 ] = 12'hf90;
    rom[1330 ] = 12'hf90;
    rom[1331 ] = 12'hf90;
    rom[1332 ] = 12'hf90;
    rom[1333 ] = 12'hf90;
    rom[1334 ] = 12'hf90;
    rom[1335 ] = 12'he90;
    rom[1336 ] = 12'he90;
    rom[1337 ] = 12'he90;
    rom[1338 ] = 12'he90;
    rom[1339 ] = 12'he90;
    rom[1340 ] = 12'he90;
    rom[1341 ] = 12'he90;
    rom[1342 ] = 12'he90;
    rom[1343 ] = 12'he90;
    rom[1344 ] = 12'he90;
    rom[1345 ] = 12'he90;
    rom[1346 ] = 12'he90;
    rom[1347 ] = 12'he90;
    rom[1348 ] = 12'he90;
    rom[1349 ] = 12'he80;
    rom[1350 ] = 12'he80;
    rom[1351 ] = 12'he80;
    rom[1352 ] = 12'he80;
    rom[1353 ] = 12'he80;
    rom[1354 ] = 12'hd80;
    rom[1355 ] = 12'hd80;
    rom[1356 ] = 12'hd80;
    rom[1357 ] = 12'hd80;
    rom[1358 ] = 12'hd80;
    rom[1359 ] = 12'hd80;
    rom[1360 ] = 12'hd80;
    rom[1361 ] = 12'hd80;
    rom[1362 ] = 12'hd80;
    rom[1363 ] = 12'hd80;
    rom[1364 ] = 12'hd80;
    rom[1365 ] = 12'hd80;
    rom[1366 ] = 12'hd80;
    rom[1367 ] = 12'hd80;
    rom[1368 ] = 12'hd80;
    rom[1369 ] = 12'hc80;
    rom[1370 ] = 12'hc80;
    rom[1371 ] = 12'hc80;
    rom[1372 ] = 12'hc80;
    rom[1373 ] = 12'hc80;
    rom[1374 ] = 12'hc80;
    rom[1375 ] = 12'hc80;
    rom[1376 ] = 12'hc80;
    rom[1377 ] = 12'hc80;
    rom[1378 ] = 12'hc80;
    rom[1379 ] = 12'h000;
    rom[1380 ] = 12'h000;
    rom[1381 ] = 12'h000;
    rom[1382 ] = 12'h000;
    rom[1383 ] = 12'h000;
    rom[1384 ] = 12'h000;
    rom[1385 ] = 12'h000;
    rom[1386 ] = 12'h000;
    rom[1387 ] = 12'h000;
    rom[1388 ] = 12'h000;
    rom[1389 ] = 12'h000;
    rom[1390 ] = 12'h000;
    rom[1391 ] = 12'h000;
    rom[1392 ] = 12'h000;
    rom[1393 ] = 12'h000;
    rom[1394 ] = 12'h000;
    rom[1395 ] = 12'h000;
    rom[1396 ] = 12'h000;
    rom[1397 ] = 12'h000;
    rom[1398 ] = 12'h000;
    rom[1399 ] = 12'h000;
    rom[1400 ] = 12'h000;
    rom[1401 ] = 12'h000;
    rom[1402 ] = 12'h000;
    rom[1403 ] = 12'h000;
    rom[1404 ] = 12'h000;
    rom[1405 ] = 12'h000;
    rom[1406 ] = 12'h000;
    rom[1407 ] = 12'h000;
    rom[1408 ] = 12'h000;
    rom[1409 ] = 12'h000;
    rom[1410 ] = 12'h000;
    rom[1411 ] = 12'h000;
    rom[1412 ] = 12'h000;
    rom[1413 ] = 12'h000;
    rom[1414 ] = 12'h000;
    rom[1415 ] = 12'h000;
    rom[1416 ] = 12'h000;
    rom[1417 ] = 12'h000;
    rom[1418 ] = 12'h000;
    rom[1419 ] = 12'h000;
    rom[1420 ] = 12'h000;
    rom[1421 ] = 12'h000;
    rom[1422 ] = 12'h000;
    rom[1423 ] = 12'h000;
    rom[1424 ] = 12'h000;
    rom[1425 ] = 12'h000;
    rom[1426 ] = 12'h000;
    rom[1427 ] = 12'h000;
    rom[1428 ] = 12'h000;
    rom[1429 ] = 12'h000;
    rom[1430 ] = 12'h000;
    rom[1431 ] = 12'h000;
    rom[1432 ] = 12'h000;
    rom[1433 ] = 12'h000;
    rom[1434 ] = 12'h000;
    rom[1435 ] = 12'h000;
    rom[1436 ] = 12'hea0;
    rom[1437 ] = 12'hea0;
    rom[1438 ] = 12'hea0;
    rom[1439 ] = 12'hea0;
    rom[1440 ] = 12'hea0;
    rom[1441 ] = 12'hea0;
    rom[1442 ] = 12'hea0;
    rom[1443 ] = 12'he90;
    rom[1444 ] = 12'hf90;
    rom[1445 ] = 12'hf90;
    rom[1446 ] = 12'hf90;
    rom[1447 ] = 12'hf90;
    rom[1448 ] = 12'hf90;
    rom[1449 ] = 12'hf90;
    rom[1450 ] = 12'hf90;
    rom[1451 ] = 12'hf90;
    rom[1452 ] = 12'hf90;
    rom[1453 ] = 12'hf90;
    rom[1454 ] = 12'hf90;
    rom[1455 ] = 12'hf90;
    rom[1456 ] = 12'hf90;
    rom[1457 ] = 12'hf90;
    rom[1458 ] = 12'hf90;
    rom[1459 ] = 12'hf90;
    rom[1460 ] = 12'hf90;
    rom[1461 ] = 12'hf90;
    rom[1462 ] = 12'hf90;
    rom[1463 ] = 12'hf90;
    rom[1464 ] = 12'he90;
    rom[1465 ] = 12'he90;
    rom[1466 ] = 12'he90;
    rom[1467 ] = 12'he90;
    rom[1468 ] = 12'he90;
    rom[1469 ] = 12'he90;
    rom[1470 ] = 12'he90;
    rom[1471 ] = 12'he90;
    rom[1472 ] = 12'he90;
    rom[1473 ] = 12'he90;
    rom[1474 ] = 12'he90;
    rom[1475 ] = 12'he90;
    rom[1476 ] = 12'he90;
    rom[1477 ] = 12'he80;
    rom[1478 ] = 12'he80;
    rom[1479 ] = 12'he80;
    rom[1480 ] = 12'he80;
    rom[1481 ] = 12'he80;
    rom[1482 ] = 12'hd80;
    rom[1483 ] = 12'hd80;
    rom[1484 ] = 12'hd80;
    rom[1485 ] = 12'hd80;
    rom[1486 ] = 12'hd80;
    rom[1487 ] = 12'hd80;
    rom[1488 ] = 12'hd80;
    rom[1489 ] = 12'hd80;
    rom[1490 ] = 12'hd80;
    rom[1491 ] = 12'hd80;
    rom[1492 ] = 12'hd80;
    rom[1493 ] = 12'hd80;
    rom[1494 ] = 12'hd80;
    rom[1495 ] = 12'hd80;
    rom[1496 ] = 12'hd80;
    rom[1497 ] = 12'hc80;
    rom[1498 ] = 12'hc80;
    rom[1499 ] = 12'hc80;
    rom[1500 ] = 12'hc80;
    rom[1501 ] = 12'hc80;
    rom[1502 ] = 12'hc80;
    rom[1503 ] = 12'hc80;
    rom[1504 ] = 12'hc80;
    rom[1505 ] = 12'hc80;
    rom[1506 ] = 12'hc80;
    rom[1507 ] = 12'hc80;
    rom[1508 ] = 12'hd90;
    rom[1509 ] = 12'h000;
    rom[1510 ] = 12'h000;
    rom[1511 ] = 12'h000;
    rom[1512 ] = 12'h000;
    rom[1513 ] = 12'h000;
    rom[1514 ] = 12'h000;
    rom[1515 ] = 12'h000;
    rom[1516 ] = 12'h000;
    rom[1517 ] = 12'h000;
    rom[1518 ] = 12'h000;
    rom[1519 ] = 12'h000;
    rom[1520 ] = 12'h000;
    rom[1521 ] = 12'h000;
    rom[1522 ] = 12'h000;
    rom[1523 ] = 12'h000;
    rom[1524 ] = 12'h000;
    rom[1525 ] = 12'h000;
    rom[1526 ] = 12'h000;
    rom[1527 ] = 12'h000;
    rom[1528 ] = 12'h000;
    rom[1529 ] = 12'h000;
    rom[1530 ] = 12'h000;
    rom[1531 ] = 12'h000;
    rom[1532 ] = 12'h000;
    rom[1533 ] = 12'h000;
    rom[1534 ] = 12'h000;
    rom[1535 ] = 12'h000;
    rom[1536 ] = 12'h000;
    rom[1537 ] = 12'h000;
    rom[1538 ] = 12'h000;
    rom[1539 ] = 12'h000;
    rom[1540 ] = 12'h000;
    rom[1541 ] = 12'h000;
    rom[1542 ] = 12'h000;
    rom[1543 ] = 12'h000;
    rom[1544 ] = 12'h000;
    rom[1545 ] = 12'h000;
    rom[1546 ] = 12'h000;
    rom[1547 ] = 12'h000;
    rom[1548 ] = 12'h000;
    rom[1549 ] = 12'h000;
    rom[1550 ] = 12'h000;
    rom[1551 ] = 12'h000;
    rom[1552 ] = 12'h000;
    rom[1553 ] = 12'h000;
    rom[1554 ] = 12'h000;
    rom[1555 ] = 12'h000;
    rom[1556 ] = 12'h000;
    rom[1557 ] = 12'h000;
    rom[1558 ] = 12'h000;
    rom[1559 ] = 12'h000;
    rom[1560 ] = 12'h000;
    rom[1561 ] = 12'h000;
    rom[1562 ] = 12'hea0;
    rom[1563 ] = 12'hea0;
    rom[1564 ] = 12'hea0;
    rom[1565 ] = 12'hea0;
    rom[1566 ] = 12'hea0;
    rom[1567 ] = 12'hea0;
    rom[1568 ] = 12'hea0;
    rom[1569 ] = 12'hea0;
    rom[1570 ] = 12'hea0;
    rom[1571 ] = 12'hea0;
    rom[1572 ] = 12'he90;
    rom[1573 ] = 12'hf90;
    rom[1574 ] = 12'hf90;
    rom[1575 ] = 12'hf90;
    rom[1576 ] = 12'hf90;
    rom[1577 ] = 12'hf90;
    rom[1578 ] = 12'hf90;
    rom[1579 ] = 12'hf90;
    rom[1580 ] = 12'hf90;
    rom[1581 ] = 12'hf90;
    rom[1582 ] = 12'hf90;
    rom[1583 ] = 12'hf90;
    rom[1584 ] = 12'hf90;
    rom[1585 ] = 12'hf90;
    rom[1586 ] = 12'hf90;
    rom[1587 ] = 12'hf90;
    rom[1588 ] = 12'hf90;
    rom[1589 ] = 12'hf90;
    rom[1590 ] = 12'hf90;
    rom[1591 ] = 12'hf90;
    rom[1592 ] = 12'he90;
    rom[1593 ] = 12'he90;
    rom[1594 ] = 12'he90;
    rom[1595 ] = 12'he90;
    rom[1596 ] = 12'he90;
    rom[1597 ] = 12'he90;
    rom[1598 ] = 12'he90;
    rom[1599 ] = 12'he90;
    rom[1600 ] = 12'he90;
    rom[1601 ] = 12'he90;
    rom[1602 ] = 12'he90;
    rom[1603 ] = 12'he90;
    rom[1604 ] = 12'he90;
    rom[1605 ] = 12'he80;
    rom[1606 ] = 12'he80;
    rom[1607 ] = 12'he80;
    rom[1608 ] = 12'he80;
    rom[1609 ] = 12'hd80;
    rom[1610 ] = 12'hd80;
    rom[1611 ] = 12'hd80;
    rom[1612 ] = 12'hd80;
    rom[1613 ] = 12'hd80;
    rom[1614 ] = 12'hd80;
    rom[1615 ] = 12'hd80;
    rom[1616 ] = 12'hd80;
    rom[1617 ] = 12'hd80;
    rom[1618 ] = 12'hd80;
    rom[1619 ] = 12'hd80;
    rom[1620 ] = 12'hd80;
    rom[1621 ] = 12'hd80;
    rom[1622 ] = 12'hd80;
    rom[1623 ] = 12'hd80;
    rom[1624 ] = 12'hc80;
    rom[1625 ] = 12'hc80;
    rom[1626 ] = 12'hc80;
    rom[1627 ] = 12'hc80;
    rom[1628 ] = 12'hc80;
    rom[1629 ] = 12'hc80;
    rom[1630 ] = 12'hc80;
    rom[1631 ] = 12'hc80;
    rom[1632 ] = 12'hc80;
    rom[1633 ] = 12'hc80;
    rom[1634 ] = 12'hc80;
    rom[1635 ] = 12'hc80;
    rom[1636 ] = 12'hc80;
    rom[1637 ] = 12'hc80;
    rom[1638 ] = 12'h000;
    rom[1639 ] = 12'h000;
    rom[1640 ] = 12'h000;
    rom[1641 ] = 12'h000;
    rom[1642 ] = 12'h000;
    rom[1643 ] = 12'h000;
    rom[1644 ] = 12'h000;
    rom[1645 ] = 12'h000;
    rom[1646 ] = 12'h000;
    rom[1647 ] = 12'h000;
    rom[1648 ] = 12'h000;
    rom[1649 ] = 12'h000;
    rom[1650 ] = 12'h000;
    rom[1651 ] = 12'h000;
    rom[1652 ] = 12'h000;
    rom[1653 ] = 12'h000;
    rom[1654 ] = 12'h000;
    rom[1655 ] = 12'h000;
    rom[1656 ] = 12'h000;
    rom[1657 ] = 12'h000;
    rom[1658 ] = 12'h000;
    rom[1659 ] = 12'h000;
    rom[1660 ] = 12'h000;
    rom[1661 ] = 12'h000;
    rom[1662 ] = 12'h000;
    rom[1663 ] = 12'h000;
    rom[1664 ] = 12'h000;
    rom[1665 ] = 12'h000;
    rom[1666 ] = 12'h000;
    rom[1667 ] = 12'h000;
    rom[1668 ] = 12'h000;
    rom[1669 ] = 12'h000;
    rom[1670 ] = 12'h000;
    rom[1671 ] = 12'h000;
    rom[1672 ] = 12'h000;
    rom[1673 ] = 12'h000;
    rom[1674 ] = 12'h000;
    rom[1675 ] = 12'h000;
    rom[1676 ] = 12'h000;
    rom[1677 ] = 12'h000;
    rom[1678 ] = 12'h000;
    rom[1679 ] = 12'h000;
    rom[1680 ] = 12'h000;
    rom[1681 ] = 12'h000;
    rom[1682 ] = 12'h000;
    rom[1683 ] = 12'h000;
    rom[1684 ] = 12'h000;
    rom[1685 ] = 12'h000;
    rom[1686 ] = 12'h000;
    rom[1687 ] = 12'h000;
    rom[1688 ] = 12'h000;
    rom[1689 ] = 12'hea0;
    rom[1690 ] = 12'hea0;
    rom[1691 ] = 12'hea0;
    rom[1692 ] = 12'hea0;
    rom[1693 ] = 12'hea0;
    rom[1694 ] = 12'hea0;
    rom[1695 ] = 12'hea0;
    rom[1696 ] = 12'hea0;
    rom[1697 ] = 12'hea0;
    rom[1698 ] = 12'hea0;
    rom[1699 ] = 12'hea0;
    rom[1700 ] = 12'he90;
    rom[1701 ] = 12'hf90;
    rom[1702 ] = 12'hf90;
    rom[1703 ] = 12'hf90;
    rom[1704 ] = 12'hf90;
    rom[1705 ] = 12'hf90;
    rom[1706 ] = 12'hf90;
    rom[1707 ] = 12'hf90;
    rom[1708 ] = 12'hf90;
    rom[1709 ] = 12'hf90;
    rom[1710 ] = 12'hf90;
    rom[1711 ] = 12'hf90;
    rom[1712 ] = 12'hf90;
    rom[1713 ] = 12'hf90;
    rom[1714 ] = 12'hf90;
    rom[1715 ] = 12'hf90;
    rom[1716 ] = 12'hf90;
    rom[1717 ] = 12'hf90;
    rom[1718 ] = 12'hf90;
    rom[1719 ] = 12'hf90;
    rom[1720 ] = 12'he90;
    rom[1721 ] = 12'he90;
    rom[1722 ] = 12'he90;
    rom[1723 ] = 12'he90;
    rom[1724 ] = 12'he90;
    rom[1725 ] = 12'he90;
    rom[1726 ] = 12'he90;
    rom[1727 ] = 12'he90;
    rom[1728 ] = 12'he90;
    rom[1729 ] = 12'he90;
    rom[1730 ] = 12'he90;
    rom[1731 ] = 12'he90;
    rom[1732 ] = 12'he80;
    rom[1733 ] = 12'he80;
    rom[1734 ] = 12'he80;
    rom[1735 ] = 12'he80;
    rom[1736 ] = 12'he80;
    rom[1737 ] = 12'hd80;
    rom[1738 ] = 12'hd80;
    rom[1739 ] = 12'hd80;
    rom[1740 ] = 12'hd80;
    rom[1741 ] = 12'hd80;
    rom[1742 ] = 12'hd80;
    rom[1743 ] = 12'hd80;
    rom[1744 ] = 12'hd80;
    rom[1745 ] = 12'hd80;
    rom[1746 ] = 12'hd80;
    rom[1747 ] = 12'hd80;
    rom[1748 ] = 12'hd80;
    rom[1749 ] = 12'hd80;
    rom[1750 ] = 12'hd80;
    rom[1751 ] = 12'hd80;
    rom[1752 ] = 12'hc80;
    rom[1753 ] = 12'hc80;
    rom[1754 ] = 12'hc80;
    rom[1755 ] = 12'hc80;
    rom[1756 ] = 12'hc80;
    rom[1757 ] = 12'hc80;
    rom[1758 ] = 12'hc80;
    rom[1759 ] = 12'hc80;
    rom[1760 ] = 12'hc80;
    rom[1761 ] = 12'hc80;
    rom[1762 ] = 12'hc80;
    rom[1763 ] = 12'hc80;
    rom[1764 ] = 12'hc80;
    rom[1765 ] = 12'hc80;
    rom[1766 ] = 12'hc80;
    rom[1767 ] = 12'h000;
    rom[1768 ] = 12'h000;
    rom[1769 ] = 12'h000;
    rom[1770 ] = 12'h000;
    rom[1771 ] = 12'h000;
    rom[1772 ] = 12'h000;
    rom[1773 ] = 12'h000;
    rom[1774 ] = 12'h000;
    rom[1775 ] = 12'h000;
    rom[1776 ] = 12'h000;
    rom[1777 ] = 12'h000;
    rom[1778 ] = 12'h000;
    rom[1779 ] = 12'h000;
    rom[1780 ] = 12'h000;
    rom[1781 ] = 12'h000;
    rom[1782 ] = 12'h000;
    rom[1783 ] = 12'h000;
    rom[1784 ] = 12'h000;
    rom[1785 ] = 12'h000;
    rom[1786 ] = 12'h000;
    rom[1787 ] = 12'h000;
    rom[1788 ] = 12'h000;
    rom[1789 ] = 12'h000;
    rom[1790 ] = 12'h000;
    rom[1791 ] = 12'h000;
    rom[1792 ] = 12'h000;
    rom[1793 ] = 12'h000;
    rom[1794 ] = 12'h000;
    rom[1795 ] = 12'h000;
    rom[1796 ] = 12'h000;
    rom[1797 ] = 12'h000;
    rom[1798 ] = 12'h000;
    rom[1799 ] = 12'h000;
    rom[1800 ] = 12'h000;
    rom[1801 ] = 12'h000;
    rom[1802 ] = 12'h000;
    rom[1803 ] = 12'h000;
    rom[1804 ] = 12'h000;
    rom[1805 ] = 12'h000;
    rom[1806 ] = 12'h000;
    rom[1807 ] = 12'h000;
    rom[1808 ] = 12'h000;
    rom[1809 ] = 12'h000;
    rom[1810 ] = 12'h000;
    rom[1811 ] = 12'h000;
    rom[1812 ] = 12'h000;
    rom[1813 ] = 12'h000;
    rom[1814 ] = 12'h000;
    rom[1815 ] = 12'h000;
    rom[1816 ] = 12'hea0;
    rom[1817 ] = 12'hea0;
    rom[1818 ] = 12'hea0;
    rom[1819 ] = 12'hea0;
    rom[1820 ] = 12'hea0;
    rom[1821 ] = 12'hea0;
    rom[1822 ] = 12'hea0;
    rom[1823 ] = 12'hea0;
    rom[1824 ] = 12'hea0;
    rom[1825 ] = 12'hea0;
    rom[1826 ] = 12'hea0;
    rom[1827 ] = 12'hea0;
    rom[1828 ] = 12'he90;
    rom[1829 ] = 12'he90;
    rom[1830 ] = 12'hf90;
    rom[1831 ] = 12'hf90;
    rom[1832 ] = 12'hf90;
    rom[1833 ] = 12'hf90;
    rom[1834 ] = 12'hf90;
    rom[1835 ] = 12'hf90;
    rom[1836 ] = 12'hf90;
    rom[1837 ] = 12'hf90;
    rom[1838 ] = 12'hf90;
    rom[1839 ] = 12'hf90;
    rom[1840 ] = 12'hf90;
    rom[1841 ] = 12'hf90;
    rom[1842 ] = 12'hf90;
    rom[1843 ] = 12'hf90;
    rom[1844 ] = 12'hf90;
    rom[1845 ] = 12'hf90;
    rom[1846 ] = 12'hf90;
    rom[1847 ] = 12'hf90;
    rom[1848 ] = 12'hf90;
    rom[1849 ] = 12'he90;
    rom[1850 ] = 12'he90;
    rom[1851 ] = 12'he90;
    rom[1852 ] = 12'he90;
    rom[1853 ] = 12'he90;
    rom[1854 ] = 12'he90;
    rom[1855 ] = 12'he90;
    rom[1856 ] = 12'he90;
    rom[1857 ] = 12'he90;
    rom[1858 ] = 12'he90;
    rom[1859 ] = 12'he90;
    rom[1860 ] = 12'he80;
    rom[1861 ] = 12'he80;
    rom[1862 ] = 12'he80;
    rom[1863 ] = 12'he80;
    rom[1864 ] = 12'he80;
    rom[1865 ] = 12'hd80;
    rom[1866 ] = 12'hd80;
    rom[1867 ] = 12'hd80;
    rom[1868 ] = 12'hd80;
    rom[1869 ] = 12'hd80;
    rom[1870 ] = 12'hd80;
    rom[1871 ] = 12'hd80;
    rom[1872 ] = 12'hd80;
    rom[1873 ] = 12'hd80;
    rom[1874 ] = 12'hd80;
    rom[1875 ] = 12'hd80;
    rom[1876 ] = 12'hd80;
    rom[1877 ] = 12'hd80;
    rom[1878 ] = 12'hd80;
    rom[1879 ] = 12'hd80;
    rom[1880 ] = 12'hc80;
    rom[1881 ] = 12'hc80;
    rom[1882 ] = 12'hc80;
    rom[1883 ] = 12'hc80;
    rom[1884 ] = 12'hc80;
    rom[1885 ] = 12'hc80;
    rom[1886 ] = 12'hc80;
    rom[1887 ] = 12'hc80;
    rom[1888 ] = 12'hc80;
    rom[1889 ] = 12'hc80;
    rom[1890 ] = 12'hc80;
    rom[1891 ] = 12'hc80;
    rom[1892 ] = 12'hc80;
    rom[1893 ] = 12'hc80;
    rom[1894 ] = 12'hc80;
    rom[1895 ] = 12'hc80;
    rom[1896 ] = 12'h000;
    rom[1897 ] = 12'h000;
    rom[1898 ] = 12'h000;
    rom[1899 ] = 12'h000;
    rom[1900 ] = 12'h000;
    rom[1901 ] = 12'h000;
    rom[1902 ] = 12'h000;
    rom[1903 ] = 12'h000;
    rom[1904 ] = 12'h000;
    rom[1905 ] = 12'h000;
    rom[1906 ] = 12'h000;
    rom[1907 ] = 12'h000;
    rom[1908 ] = 12'h000;
    rom[1909 ] = 12'h000;
    rom[1910 ] = 12'h000;
    rom[1911 ] = 12'h000;
    rom[1912 ] = 12'h000;
    rom[1913 ] = 12'h000;
    rom[1914 ] = 12'h000;
    rom[1915 ] = 12'h000;
    rom[1916 ] = 12'h000;
    rom[1917 ] = 12'h000;
    rom[1918 ] = 12'h000;
    rom[1919 ] = 12'h000;
    rom[1920 ] = 12'h000;
    rom[1921 ] = 12'h000;
    rom[1922 ] = 12'h000;
    rom[1923 ] = 12'h000;
    rom[1924 ] = 12'h000;
    rom[1925 ] = 12'h000;
    rom[1926 ] = 12'h000;
    rom[1927 ] = 12'h000;
    rom[1928 ] = 12'h000;
    rom[1929 ] = 12'h000;
    rom[1930 ] = 12'h000;
    rom[1931 ] = 12'h000;
    rom[1932 ] = 12'h000;
    rom[1933 ] = 12'h000;
    rom[1934 ] = 12'h000;
    rom[1935 ] = 12'h000;
    rom[1936 ] = 12'h000;
    rom[1937 ] = 12'h000;
    rom[1938 ] = 12'h000;
    rom[1939 ] = 12'h000;
    rom[1940 ] = 12'h000;
    rom[1941 ] = 12'h000;
    rom[1942 ] = 12'hda0;
    rom[1943 ] = 12'hea0;
    rom[1944 ] = 12'hea0;
    rom[1945 ] = 12'hea0;
    rom[1946 ] = 12'hea0;
    rom[1947 ] = 12'hea0;
    rom[1948 ] = 12'hea0;
    rom[1949 ] = 12'hea0;
    rom[1950 ] = 12'hea0;
    rom[1951 ] = 12'hea0;
    rom[1952 ] = 12'hea0;
    rom[1953 ] = 12'hea0;
    rom[1954 ] = 12'hea0;
    rom[1955 ] = 12'hea0;
    rom[1956 ] = 12'hea0;
    rom[1957 ] = 12'he90;
    rom[1958 ] = 12'hf90;
    rom[1959 ] = 12'hf90;
    rom[1960 ] = 12'hf90;
    rom[1961 ] = 12'hf90;
    rom[1962 ] = 12'hf90;
    rom[1963 ] = 12'hf90;
    rom[1964 ] = 12'hf90;
    rom[1965 ] = 12'hf90;
    rom[1966 ] = 12'hf90;
    rom[1967 ] = 12'hf90;
    rom[1968 ] = 12'hf90;
    rom[1969 ] = 12'hf90;
    rom[1970 ] = 12'hf90;
    rom[1971 ] = 12'hf90;
    rom[1972 ] = 12'hf90;
    rom[1973 ] = 12'hf90;
    rom[1974 ] = 12'hf90;
    rom[1975 ] = 12'hf90;
    rom[1976 ] = 12'hf90;
    rom[1977 ] = 12'h000;
    rom[1978 ] = 12'h000;
    rom[1979 ] = 12'h000;
    rom[1980 ] = 12'h000;
    rom[1981 ] = 12'h000;
    rom[1982 ] = 12'h000;
    rom[1983 ] = 12'h000;
    rom[1984 ] = 12'h000;
    rom[1985 ] = 12'h000;
    rom[1986 ] = 12'h000;
    rom[1987 ] = 12'h000;
    rom[1988 ] = 12'h000;
    rom[1989 ] = 12'h000;
    rom[1990 ] = 12'h000;
    rom[1991 ] = 12'he80;
    rom[1992 ] = 12'hd80;
    rom[1993 ] = 12'hd80;
    rom[1994 ] = 12'hd80;
    rom[1995 ] = 12'hd80;
    rom[1996 ] = 12'hd80;
    rom[1997 ] = 12'hd80;
    rom[1998 ] = 12'hd80;
    rom[1999 ] = 12'hd80;
    rom[2000 ] = 12'hd80;
    rom[2001 ] = 12'hd80;
    rom[2002 ] = 12'hd80;
    rom[2003 ] = 12'hd80;
    rom[2004 ] = 12'hd80;
    rom[2005 ] = 12'hd80;
    rom[2006 ] = 12'hd80;
    rom[2007 ] = 12'hd80;
    rom[2008 ] = 12'hc80;
    rom[2009 ] = 12'hc80;
    rom[2010 ] = 12'hc80;
    rom[2011 ] = 12'hc80;
    rom[2012 ] = 12'hc80;
    rom[2013 ] = 12'hc80;
    rom[2014 ] = 12'hc80;
    rom[2015 ] = 12'hc80;
    rom[2016 ] = 12'hc80;
    rom[2017 ] = 12'hc80;
    rom[2018 ] = 12'hc80;
    rom[2019 ] = 12'hc80;
    rom[2020 ] = 12'hc80;
    rom[2021 ] = 12'hc80;
    rom[2022 ] = 12'hc80;
    rom[2023 ] = 12'h000;
    rom[2024 ] = 12'h000;
    rom[2025 ] = 12'h000;
    rom[2026 ] = 12'h000;
    rom[2027 ] = 12'h000;
    rom[2028 ] = 12'h000;
    rom[2029 ] = 12'h000;
    rom[2030 ] = 12'h000;
    rom[2031 ] = 12'h000;
    rom[2032 ] = 12'h000;
    rom[2033 ] = 12'h000;
    rom[2034 ] = 12'h000;
    rom[2035 ] = 12'h000;
    rom[2036 ] = 12'h000;
    rom[2037 ] = 12'h000;
    rom[2038 ] = 12'h000;
    rom[2039 ] = 12'h000;
    rom[2040 ] = 12'h000;
    rom[2041 ] = 12'h000;
    rom[2042 ] = 12'h000;
    rom[2043 ] = 12'h000;
    rom[2044 ] = 12'h000;
    rom[2045 ] = 12'h000;
    rom[2046 ] = 12'h000;
    rom[2047 ] = 12'h000;
    rom[2048 ] = 12'h000;
    rom[2049 ] = 12'h000;
    rom[2050 ] = 12'h000;
    rom[2051 ] = 12'h000;
    rom[2052 ] = 12'h000;
    rom[2053 ] = 12'h000;
    rom[2054 ] = 12'h000;
    rom[2055 ] = 12'h000;
    rom[2056 ] = 12'h000;
    rom[2057 ] = 12'h000;
    rom[2058 ] = 12'h000;
    rom[2059 ] = 12'h000;
    rom[2060 ] = 12'h000;
    rom[2061 ] = 12'h000;
    rom[2062 ] = 12'h000;
    rom[2063 ] = 12'h000;
    rom[2064 ] = 12'h000;
    rom[2065 ] = 12'h000;
    rom[2066 ] = 12'h000;
    rom[2067 ] = 12'h000;
    rom[2068 ] = 12'h000;
    rom[2069 ] = 12'hea0;
    rom[2070 ] = 12'hea0;
    rom[2071 ] = 12'hea0;
    rom[2072 ] = 12'hea0;
    rom[2073 ] = 12'hea0;
    rom[2074 ] = 12'hea0;
    rom[2075 ] = 12'hea0;
    rom[2076 ] = 12'hea0;
    rom[2077 ] = 12'hea0;
    rom[2078 ] = 12'hea0;
    rom[2079 ] = 12'hea0;
    rom[2080 ] = 12'hea0;
    rom[2081 ] = 12'hea0;
    rom[2082 ] = 12'hea0;
    rom[2083 ] = 12'hea0;
    rom[2084 ] = 12'hea0;
    rom[2085 ] = 12'he90;
    rom[2086 ] = 12'hf90;
    rom[2087 ] = 12'hf90;
    rom[2088 ] = 12'hf90;
    rom[2089 ] = 12'hf90;
    rom[2090 ] = 12'hf90;
    rom[2091 ] = 12'hf90;
    rom[2092 ] = 12'hf90;
    rom[2093 ] = 12'hf90;
    rom[2094 ] = 12'hf90;
    rom[2095 ] = 12'hf90;
    rom[2096 ] = 12'hf90;
    rom[2097 ] = 12'hf90;
    rom[2098 ] = 12'hf90;
    rom[2099 ] = 12'hf90;
    rom[2100 ] = 12'h000;
    rom[2101 ] = 12'h000;
    rom[2102 ] = 12'h000;
    rom[2103 ] = 12'h000;
    rom[2104 ] = 12'h000;
    rom[2105 ] = 12'h000;
    rom[2106 ] = 12'h000;
    rom[2107 ] = 12'h000;
    rom[2108 ] = 12'h000;
    rom[2109 ] = 12'h000;
    rom[2110 ] = 12'h000;
    rom[2111 ] = 12'h000;
    rom[2112 ] = 12'h000;
    rom[2113 ] = 12'h000;
    rom[2114 ] = 12'h000;
    rom[2115 ] = 12'h000;
    rom[2116 ] = 12'h000;
    rom[2117 ] = 12'h000;
    rom[2118 ] = 12'h000;
    rom[2119 ] = 12'h000;
    rom[2120 ] = 12'h000;
    rom[2121 ] = 12'h000;
    rom[2122 ] = 12'h000;
    rom[2123 ] = 12'h000;
    rom[2124 ] = 12'hd80;
    rom[2125 ] = 12'hd80;
    rom[2126 ] = 12'hd80;
    rom[2127 ] = 12'hd80;
    rom[2128 ] = 12'hd80;
    rom[2129 ] = 12'hd80;
    rom[2130 ] = 12'hd80;
    rom[2131 ] = 12'hd80;
    rom[2132 ] = 12'hd80;
    rom[2133 ] = 12'hd80;
    rom[2134 ] = 12'hd80;
    rom[2135 ] = 12'hc80;
    rom[2136 ] = 12'hc80;
    rom[2137 ] = 12'hc80;
    rom[2138 ] = 12'hc80;
    rom[2139 ] = 12'hc80;
    rom[2140 ] = 12'hc80;
    rom[2141 ] = 12'hc80;
    rom[2142 ] = 12'hc80;
    rom[2143 ] = 12'hc80;
    rom[2144 ] = 12'hc80;
    rom[2145 ] = 12'hc80;
    rom[2146 ] = 12'hc80;
    rom[2147 ] = 12'hc80;
    rom[2148 ] = 12'hc80;
    rom[2149 ] = 12'h000;
    rom[2150 ] = 12'h000;
    rom[2151 ] = 12'h000;
    rom[2152 ] = 12'h000;
    rom[2153 ] = 12'h000;
    rom[2154 ] = 12'h000;
    rom[2155 ] = 12'h000;
    rom[2156 ] = 12'h000;
    rom[2157 ] = 12'h000;
    rom[2158 ] = 12'h000;
    rom[2159 ] = 12'h000;
    rom[2160 ] = 12'h000;
    rom[2161 ] = 12'h000;
    rom[2162 ] = 12'h000;
    rom[2163 ] = 12'h000;
    rom[2164 ] = 12'h000;
    rom[2165 ] = 12'h000;
    rom[2166 ] = 12'h000;
    rom[2167 ] = 12'h000;
    rom[2168 ] = 12'h000;
    rom[2169 ] = 12'h000;
    rom[2170 ] = 12'h000;
    rom[2171 ] = 12'h000;
    rom[2172 ] = 12'h000;
    rom[2173 ] = 12'h000;
    rom[2174 ] = 12'h000;
    rom[2175 ] = 12'h000;
    rom[2176 ] = 12'h000;
    rom[2177 ] = 12'h000;
    rom[2178 ] = 12'h000;
    rom[2179 ] = 12'h000;
    rom[2180 ] = 12'h000;
    rom[2181 ] = 12'h000;
    rom[2182 ] = 12'h000;
    rom[2183 ] = 12'h000;
    rom[2184 ] = 12'h000;
    rom[2185 ] = 12'h000;
    rom[2186 ] = 12'h000;
    rom[2187 ] = 12'h000;
    rom[2188 ] = 12'h000;
    rom[2189 ] = 12'h000;
    rom[2190 ] = 12'h000;
    rom[2191 ] = 12'h000;
    rom[2192 ] = 12'h000;
    rom[2193 ] = 12'h000;
    rom[2194 ] = 12'h000;
    rom[2195 ] = 12'h000;
    rom[2196 ] = 12'hea0;
    rom[2197 ] = 12'hea0;
    rom[2198 ] = 12'hea0;
    rom[2199 ] = 12'hea0;
    rom[2200 ] = 12'hea0;
    rom[2201 ] = 12'hea0;
    rom[2202 ] = 12'hea0;
    rom[2203 ] = 12'hea0;
    rom[2204 ] = 12'hea0;
    rom[2205 ] = 12'hea0;
    rom[2206 ] = 12'hea0;
    rom[2207 ] = 12'hea0;
    rom[2208 ] = 12'hea0;
    rom[2209 ] = 12'hea0;
    rom[2210 ] = 12'hea0;
    rom[2211 ] = 12'hea0;
    rom[2212 ] = 12'hea0;
    rom[2213 ] = 12'hea0;
    rom[2214 ] = 12'he90;
    rom[2215 ] = 12'hf90;
    rom[2216 ] = 12'hf90;
    rom[2217 ] = 12'hf90;
    rom[2218 ] = 12'hf90;
    rom[2219 ] = 12'hf90;
    rom[2220 ] = 12'hf90;
    rom[2221 ] = 12'hf90;
    rom[2222 ] = 12'hf90;
    rom[2223 ] = 12'hf90;
    rom[2224 ] = 12'hf90;
    rom[2225 ] = 12'h000;
    rom[2226 ] = 12'h000;
    rom[2227 ] = 12'h000;
    rom[2228 ] = 12'h000;
    rom[2229 ] = 12'h000;
    rom[2230 ] = 12'h000;
    rom[2231 ] = 12'h000;
    rom[2232 ] = 12'h000;
    rom[2233 ] = 12'h000;
    rom[2234 ] = 12'h000;
    rom[2235 ] = 12'h000;
    rom[2236 ] = 12'h000;
    rom[2237 ] = 12'h000;
    rom[2238 ] = 12'h000;
    rom[2239 ] = 12'h000;
    rom[2240 ] = 12'h000;
    rom[2241 ] = 12'h000;
    rom[2242 ] = 12'h000;
    rom[2243 ] = 12'h000;
    rom[2244 ] = 12'h000;
    rom[2245 ] = 12'h000;
    rom[2246 ] = 12'h000;
    rom[2247 ] = 12'h000;
    rom[2248 ] = 12'h000;
    rom[2249 ] = 12'h000;
    rom[2250 ] = 12'h000;
    rom[2251 ] = 12'h000;
    rom[2252 ] = 12'h000;
    rom[2253 ] = 12'h000;
    rom[2254 ] = 12'h000;
    rom[2255 ] = 12'hd80;
    rom[2256 ] = 12'hd80;
    rom[2257 ] = 12'hd80;
    rom[2258 ] = 12'hd80;
    rom[2259 ] = 12'hd80;
    rom[2260 ] = 12'hd80;
    rom[2261 ] = 12'hd80;
    rom[2262 ] = 12'hd80;
    rom[2263 ] = 12'hc80;
    rom[2264 ] = 12'hc80;
    rom[2265 ] = 12'hc80;
    rom[2266 ] = 12'hc80;
    rom[2267 ] = 12'hc80;
    rom[2268 ] = 12'hc80;
    rom[2269 ] = 12'hc80;
    rom[2270 ] = 12'hc80;
    rom[2271 ] = 12'hc80;
    rom[2272 ] = 12'hc80;
    rom[2273 ] = 12'hc80;
    rom[2274 ] = 12'hc80;
    rom[2275 ] = 12'hc80;
    rom[2276 ] = 12'h000;
    rom[2277 ] = 12'h000;
    rom[2278 ] = 12'h000;
    rom[2279 ] = 12'h000;
    rom[2280 ] = 12'h000;
    rom[2281 ] = 12'h000;
    rom[2282 ] = 12'h000;
    rom[2283 ] = 12'h000;
    rom[2284 ] = 12'h000;
    rom[2285 ] = 12'h000;
    rom[2286 ] = 12'h000;
    rom[2287 ] = 12'h000;
    rom[2288 ] = 12'h000;
    rom[2289 ] = 12'h000;
    rom[2290 ] = 12'h000;
    rom[2291 ] = 12'h000;
    rom[2292 ] = 12'h000;
    rom[2293 ] = 12'h000;
    rom[2294 ] = 12'h000;
    rom[2295 ] = 12'h000;
    rom[2296 ] = 12'h000;
    rom[2297 ] = 12'h000;
    rom[2298 ] = 12'h000;
    rom[2299 ] = 12'h000;
    rom[2300 ] = 12'h000;
    rom[2301 ] = 12'h000;
    rom[2302 ] = 12'h000;
    rom[2303 ] = 12'h000;
    rom[2304 ] = 12'h000;
    rom[2305 ] = 12'h000;
    rom[2306 ] = 12'h000;
    rom[2307 ] = 12'h000;
    rom[2308 ] = 12'h000;
    rom[2309 ] = 12'h000;
    rom[2310 ] = 12'h000;
    rom[2311 ] = 12'h000;
    rom[2312 ] = 12'h000;
    rom[2313 ] = 12'h000;
    rom[2314 ] = 12'h000;
    rom[2315 ] = 12'h000;
    rom[2316 ] = 12'h000;
    rom[2317 ] = 12'h000;
    rom[2318 ] = 12'h000;
    rom[2319 ] = 12'h000;
    rom[2320 ] = 12'h000;
    rom[2321 ] = 12'h000;
    rom[2322 ] = 12'h000;
    rom[2323 ] = 12'hea0;
    rom[2324 ] = 12'hea0;
    rom[2325 ] = 12'hea0;
    rom[2326 ] = 12'hea0;
    rom[2327 ] = 12'hea0;
    rom[2328 ] = 12'hea0;
    rom[2329 ] = 12'hea0;
    rom[2330 ] = 12'hea0;
    rom[2331 ] = 12'hea0;
    rom[2332 ] = 12'hea0;
    rom[2333 ] = 12'hea0;
    rom[2334 ] = 12'hea0;
    rom[2335 ] = 12'hea0;
    rom[2336 ] = 12'hea0;
    rom[2337 ] = 12'hea0;
    rom[2338 ] = 12'hea0;
    rom[2339 ] = 12'hea0;
    rom[2340 ] = 12'hea0;
    rom[2341 ] = 12'hea0;
    rom[2342 ] = 12'he90;
    rom[2343 ] = 12'hf90;
    rom[2344 ] = 12'hf90;
    rom[2345 ] = 12'hf90;
    rom[2346 ] = 12'hf90;
    rom[2347 ] = 12'hf90;
    rom[2348 ] = 12'hf90;
    rom[2349 ] = 12'hf90;
    rom[2350 ] = 12'h000;
    rom[2351 ] = 12'h000;
    rom[2352 ] = 12'h000;
    rom[2353 ] = 12'h000;
    rom[2354 ] = 12'h000;
    rom[2355 ] = 12'h000;
    rom[2356 ] = 12'h000;
    rom[2357 ] = 12'h000;
    rom[2358 ] = 12'h000;
    rom[2359 ] = 12'h000;
    rom[2360 ] = 12'h000;
    rom[2361 ] = 12'h000;
    rom[2362 ] = 12'h000;
    rom[2363 ] = 12'h000;
    rom[2364 ] = 12'h000;
    rom[2365 ] = 12'h000;
    rom[2366 ] = 12'h000;
    rom[2367 ] = 12'h000;
    rom[2368 ] = 12'h000;
    rom[2369 ] = 12'h000;
    rom[2370 ] = 12'h000;
    rom[2371 ] = 12'h000;
    rom[2372 ] = 12'h000;
    rom[2373 ] = 12'h000;
    rom[2374 ] = 12'h000;
    rom[2375 ] = 12'h000;
    rom[2376 ] = 12'h000;
    rom[2377 ] = 12'h000;
    rom[2378 ] = 12'h000;
    rom[2379 ] = 12'h000;
    rom[2380 ] = 12'h000;
    rom[2381 ] = 12'h000;
    rom[2382 ] = 12'h000;
    rom[2383 ] = 12'h000;
    rom[2384 ] = 12'h000;
    rom[2385 ] = 12'h000;
    rom[2386 ] = 12'hd80;
    rom[2387 ] = 12'hd80;
    rom[2388 ] = 12'hd80;
    rom[2389 ] = 12'hd80;
    rom[2390 ] = 12'hd80;
    rom[2391 ] = 12'hc80;
    rom[2392 ] = 12'hc80;
    rom[2393 ] = 12'hc80;
    rom[2394 ] = 12'hc80;
    rom[2395 ] = 12'hc80;
    rom[2396 ] = 12'hc80;
    rom[2397 ] = 12'hc80;
    rom[2398 ] = 12'hc80;
    rom[2399 ] = 12'hc80;
    rom[2400 ] = 12'hc80;
    rom[2401 ] = 12'hc80;
    rom[2402 ] = 12'hc80;
    rom[2403 ] = 12'h000;
    rom[2404 ] = 12'h000;
    rom[2405 ] = 12'h000;
    rom[2406 ] = 12'h000;
    rom[2407 ] = 12'h000;
    rom[2408 ] = 12'h000;
    rom[2409 ] = 12'h000;
    rom[2410 ] = 12'h000;
    rom[2411 ] = 12'h000;
    rom[2412 ] = 12'h000;
    rom[2413 ] = 12'h000;
    rom[2414 ] = 12'h000;
    rom[2415 ] = 12'h000;
    rom[2416 ] = 12'h000;
    rom[2417 ] = 12'h000;
    rom[2418 ] = 12'h000;
    rom[2419 ] = 12'h000;
    rom[2420 ] = 12'h000;
    rom[2421 ] = 12'h000;
    rom[2422 ] = 12'h000;
    rom[2423 ] = 12'h000;
    rom[2424 ] = 12'h000;
    rom[2425 ] = 12'h000;
    rom[2426 ] = 12'h000;
    rom[2427 ] = 12'h000;
    rom[2428 ] = 12'h000;
    rom[2429 ] = 12'h000;
    rom[2430 ] = 12'h000;
    rom[2431 ] = 12'h000;
    rom[2432 ] = 12'h000;
    rom[2433 ] = 12'h000;
    rom[2434 ] = 12'h000;
    rom[2435 ] = 12'h000;
    rom[2436 ] = 12'h000;
    rom[2437 ] = 12'h000;
    rom[2438 ] = 12'h000;
    rom[2439 ] = 12'h000;
    rom[2440 ] = 12'h000;
    rom[2441 ] = 12'h000;
    rom[2442 ] = 12'h000;
    rom[2443 ] = 12'h000;
    rom[2444 ] = 12'h000;
    rom[2445 ] = 12'h000;
    rom[2446 ] = 12'h000;
    rom[2447 ] = 12'h000;
    rom[2448 ] = 12'h000;
    rom[2449 ] = 12'h000;
    rom[2450 ] = 12'hea0;
    rom[2451 ] = 12'hea0;
    rom[2452 ] = 12'hea0;
    rom[2453 ] = 12'hea0;
    rom[2454 ] = 12'hea0;
    rom[2455 ] = 12'hea0;
    rom[2456 ] = 12'hea0;
    rom[2457 ] = 12'hea0;
    rom[2458 ] = 12'hea0;
    rom[2459 ] = 12'hea0;
    rom[2460 ] = 12'hea0;
    rom[2461 ] = 12'hea0;
    rom[2462 ] = 12'hea0;
    rom[2463 ] = 12'hea0;
    rom[2464 ] = 12'hea0;
    rom[2465 ] = 12'hea0;
    rom[2466 ] = 12'hea0;
    rom[2467 ] = 12'hea0;
    rom[2468 ] = 12'hea0;
    rom[2469 ] = 12'hea0;
    rom[2470 ] = 12'he90;
    rom[2471 ] = 12'hf90;
    rom[2472 ] = 12'hf90;
    rom[2473 ] = 12'hf90;
    rom[2474 ] = 12'hf90;
    rom[2475 ] = 12'hfa0;
    rom[2476 ] = 12'h000;
    rom[2477 ] = 12'h000;
    rom[2478 ] = 12'h000;
    rom[2479 ] = 12'h000;
    rom[2480 ] = 12'h000;
    rom[2481 ] = 12'h000;
    rom[2482 ] = 12'h000;
    rom[2483 ] = 12'h000;
    rom[2484 ] = 12'h000;
    rom[2485 ] = 12'h000;
    rom[2486 ] = 12'h000;
    rom[2487 ] = 12'h000;
    rom[2488 ] = 12'h000;
    rom[2489 ] = 12'h000;
    rom[2490 ] = 12'h000;
    rom[2491 ] = 12'h000;
    rom[2492 ] = 12'h000;
    rom[2493 ] = 12'h000;
    rom[2494 ] = 12'h000;
    rom[2495 ] = 12'h000;
    rom[2496 ] = 12'h000;
    rom[2497 ] = 12'h000;
    rom[2498 ] = 12'h000;
    rom[2499 ] = 12'h000;
    rom[2500 ] = 12'h000;
    rom[2501 ] = 12'h000;
    rom[2502 ] = 12'h000;
    rom[2503 ] = 12'h000;
    rom[2504 ] = 12'h000;
    rom[2505 ] = 12'h000;
    rom[2506 ] = 12'h000;
    rom[2507 ] = 12'h000;
    rom[2508 ] = 12'h000;
    rom[2509 ] = 12'h000;
    rom[2510 ] = 12'h000;
    rom[2511 ] = 12'h000;
    rom[2512 ] = 12'h000;
    rom[2513 ] = 12'h000;
    rom[2514 ] = 12'h000;
    rom[2515 ] = 12'h000;
    rom[2516 ] = 12'hd80;
    rom[2517 ] = 12'hd80;
    rom[2518 ] = 12'hc80;
    rom[2519 ] = 12'hc80;
    rom[2520 ] = 12'hc80;
    rom[2521 ] = 12'hc80;
    rom[2522 ] = 12'hc80;
    rom[2523 ] = 12'hc80;
    rom[2524 ] = 12'hc80;
    rom[2525 ] = 12'hc80;
    rom[2526 ] = 12'hc80;
    rom[2527 ] = 12'hc80;
    rom[2528 ] = 12'hc80;
    rom[2529 ] = 12'h000;
    rom[2530 ] = 12'h000;
    rom[2531 ] = 12'h000;
    rom[2532 ] = 12'h000;
    rom[2533 ] = 12'h000;
    rom[2534 ] = 12'h000;
    rom[2535 ] = 12'h000;
    rom[2536 ] = 12'h000;
    rom[2537 ] = 12'h000;
    rom[2538 ] = 12'h000;
    rom[2539 ] = 12'h000;
    rom[2540 ] = 12'h000;
    rom[2541 ] = 12'h000;
    rom[2542 ] = 12'h000;
    rom[2543 ] = 12'h000;
    rom[2544 ] = 12'h000;
    rom[2545 ] = 12'h000;
    rom[2546 ] = 12'h000;
    rom[2547 ] = 12'h000;
    rom[2548 ] = 12'h000;
    rom[2549 ] = 12'h000;
    rom[2550 ] = 12'h000;
    rom[2551 ] = 12'h000;
    rom[2552 ] = 12'h000;
    rom[2553 ] = 12'h000;
    rom[2554 ] = 12'h000;
    rom[2555 ] = 12'h000;
    rom[2556 ] = 12'h000;
    rom[2557 ] = 12'h000;
    rom[2558 ] = 12'h000;
    rom[2559 ] = 12'h000;
    rom[2560 ] = 12'h000;
    rom[2561 ] = 12'h000;
    rom[2562 ] = 12'h000;
    rom[2563 ] = 12'h000;
    rom[2564 ] = 12'h000;
    rom[2565 ] = 12'h000;
    rom[2566 ] = 12'h000;
    rom[2567 ] = 12'h000;
    rom[2568 ] = 12'h000;
    rom[2569 ] = 12'h000;
    rom[2570 ] = 12'h000;
    rom[2571 ] = 12'h000;
    rom[2572 ] = 12'h000;
    rom[2573 ] = 12'h000;
    rom[2574 ] = 12'h000;
    rom[2575 ] = 12'h000;
    rom[2576 ] = 12'h000;
    rom[2577 ] = 12'hea0;
    rom[2578 ] = 12'hea0;
    rom[2579 ] = 12'hea0;
    rom[2580 ] = 12'hea0;
    rom[2581 ] = 12'hea0;
    rom[2582 ] = 12'hea0;
    rom[2583 ] = 12'hea0;
    rom[2584 ] = 12'hea0;
    rom[2585 ] = 12'hea0;
    rom[2586 ] = 12'hea0;
    rom[2587 ] = 12'hea0;
    rom[2588 ] = 12'hea0;
    rom[2589 ] = 12'hea0;
    rom[2590 ] = 12'hea0;
    rom[2591 ] = 12'hea0;
    rom[2592 ] = 12'hea0;
    rom[2593 ] = 12'hea0;
    rom[2594 ] = 12'hea0;
    rom[2595 ] = 12'hea0;
    rom[2596 ] = 12'hea0;
    rom[2597 ] = 12'hea0;
    rom[2598 ] = 12'hea0;
    rom[2599 ] = 12'he90;
    rom[2600 ] = 12'hf90;
    rom[2601 ] = 12'hf90;
    rom[2602 ] = 12'h000;
    rom[2603 ] = 12'h000;
    rom[2604 ] = 12'h000;
    rom[2605 ] = 12'h000;
    rom[2606 ] = 12'h000;
    rom[2607 ] = 12'h000;
    rom[2608 ] = 12'h000;
    rom[2609 ] = 12'h000;
    rom[2610 ] = 12'h000;
    rom[2611 ] = 12'h000;
    rom[2612 ] = 12'h000;
    rom[2613 ] = 12'h000;
    rom[2614 ] = 12'h000;
    rom[2615 ] = 12'h000;
    rom[2616 ] = 12'h000;
    rom[2617 ] = 12'h000;
    rom[2618 ] = 12'h000;
    rom[2619 ] = 12'h000;
    rom[2620 ] = 12'h000;
    rom[2621 ] = 12'h000;
    rom[2622 ] = 12'h000;
    rom[2623 ] = 12'h000;
    rom[2624 ] = 12'h000;
    rom[2625 ] = 12'h000;
    rom[2626 ] = 12'h000;
    rom[2627 ] = 12'h000;
    rom[2628 ] = 12'h000;
    rom[2629 ] = 12'h000;
    rom[2630 ] = 12'h000;
    rom[2631 ] = 12'h000;
    rom[2632 ] = 12'h000;
    rom[2633 ] = 12'h000;
    rom[2634 ] = 12'h000;
    rom[2635 ] = 12'h000;
    rom[2636 ] = 12'h000;
    rom[2637 ] = 12'h000;
    rom[2638 ] = 12'h000;
    rom[2639 ] = 12'h000;
    rom[2640 ] = 12'h000;
    rom[2641 ] = 12'h000;
    rom[2642 ] = 12'h000;
    rom[2643 ] = 12'h000;
    rom[2644 ] = 12'h000;
    rom[2645 ] = 12'h000;
    rom[2646 ] = 12'hd91;
    rom[2647 ] = 12'hc80;
    rom[2648 ] = 12'hc80;
    rom[2649 ] = 12'hc80;
    rom[2650 ] = 12'hc80;
    rom[2651 ] = 12'hc80;
    rom[2652 ] = 12'hc80;
    rom[2653 ] = 12'hc80;
    rom[2654 ] = 12'hc80;
    rom[2655 ] = 12'hc80;
    rom[2656 ] = 12'h000;
    rom[2657 ] = 12'h000;
    rom[2658 ] = 12'h000;
    rom[2659 ] = 12'h000;
    rom[2660 ] = 12'h000;
    rom[2661 ] = 12'h000;
    rom[2662 ] = 12'h000;
    rom[2663 ] = 12'h000;
    rom[2664 ] = 12'h000;
    rom[2665 ] = 12'h000;
    rom[2666 ] = 12'h000;
    rom[2667 ] = 12'h000;
    rom[2668 ] = 12'h000;
    rom[2669 ] = 12'h000;
    rom[2670 ] = 12'h000;
    rom[2671 ] = 12'h000;
    rom[2672 ] = 12'h000;
    rom[2673 ] = 12'h000;
    rom[2674 ] = 12'h000;
    rom[2675 ] = 12'h000;
    rom[2676 ] = 12'h000;
    rom[2677 ] = 12'h000;
    rom[2678 ] = 12'h000;
    rom[2679 ] = 12'h000;
    rom[2680 ] = 12'h000;
    rom[2681 ] = 12'h000;
    rom[2682 ] = 12'h000;
    rom[2683 ] = 12'h000;
    rom[2684 ] = 12'h000;
    rom[2685 ] = 12'h000;
    rom[2686 ] = 12'h000;
    rom[2687 ] = 12'h000;
    rom[2688 ] = 12'h000;
    rom[2689 ] = 12'h000;
    rom[2690 ] = 12'h000;
    rom[2691 ] = 12'h000;
    rom[2692 ] = 12'h000;
    rom[2693 ] = 12'h000;
    rom[2694 ] = 12'h000;
    rom[2695 ] = 12'h000;
    rom[2696 ] = 12'h000;
    rom[2697 ] = 12'h000;
    rom[2698 ] = 12'h000;
    rom[2699 ] = 12'h000;
    rom[2700 ] = 12'h000;
    rom[2701 ] = 12'h000;
    rom[2702 ] = 12'h000;
    rom[2703 ] = 12'h000;
    rom[2704 ] = 12'hea0;
    rom[2705 ] = 12'hea0;
    rom[2706 ] = 12'hea0;
    rom[2707 ] = 12'hea0;
    rom[2708 ] = 12'hea0;
    rom[2709 ] = 12'hea0;
    rom[2710 ] = 12'hea0;
    rom[2711 ] = 12'hea0;
    rom[2712 ] = 12'hea0;
    rom[2713 ] = 12'hea0;
    rom[2714 ] = 12'hea0;
    rom[2715 ] = 12'hea0;
    rom[2716 ] = 12'hea0;
    rom[2717 ] = 12'hea0;
    rom[2718 ] = 12'hea0;
    rom[2719 ] = 12'hea0;
    rom[2720 ] = 12'hea0;
    rom[2721 ] = 12'hea0;
    rom[2722 ] = 12'hea0;
    rom[2723 ] = 12'hea0;
    rom[2724 ] = 12'hea0;
    rom[2725 ] = 12'hea0;
    rom[2726 ] = 12'hea0;
    rom[2727 ] = 12'he90;
    rom[2728 ] = 12'h000;
    rom[2729 ] = 12'h000;
    rom[2730 ] = 12'h000;
    rom[2731 ] = 12'h000;
    rom[2732 ] = 12'h000;
    rom[2733 ] = 12'h000;
    rom[2734 ] = 12'h000;
    rom[2735 ] = 12'h000;
    rom[2736 ] = 12'h000;
    rom[2737 ] = 12'h000;
    rom[2738 ] = 12'h000;
    rom[2739 ] = 12'h000;
    rom[2740 ] = 12'h000;
    rom[2741 ] = 12'h000;
    rom[2742 ] = 12'h000;
    rom[2743 ] = 12'h000;
    rom[2744 ] = 12'h000;
    rom[2745 ] = 12'h000;
    rom[2746 ] = 12'h000;
    rom[2747 ] = 12'h000;
    rom[2748 ] = 12'h000;
    rom[2749 ] = 12'h000;
    rom[2750 ] = 12'h000;
    rom[2751 ] = 12'h000;
    rom[2752 ] = 12'h000;
    rom[2753 ] = 12'h000;
    rom[2754 ] = 12'h000;
    rom[2755 ] = 12'h000;
    rom[2756 ] = 12'h000;
    rom[2757 ] = 12'h000;
    rom[2758 ] = 12'h000;
    rom[2759 ] = 12'h000;
    rom[2760 ] = 12'h000;
    rom[2761 ] = 12'h000;
    rom[2762 ] = 12'h000;
    rom[2763 ] = 12'h000;
    rom[2764 ] = 12'h000;
    rom[2765 ] = 12'h000;
    rom[2766 ] = 12'h000;
    rom[2767 ] = 12'h000;
    rom[2768 ] = 12'h000;
    rom[2769 ] = 12'h000;
    rom[2770 ] = 12'h000;
    rom[2771 ] = 12'h000;
    rom[2772 ] = 12'h000;
    rom[2773 ] = 12'h000;
    rom[2774 ] = 12'h000;
    rom[2775 ] = 12'h000;
    rom[2776 ] = 12'hc80;
    rom[2777 ] = 12'hc80;
    rom[2778 ] = 12'hc80;
    rom[2779 ] = 12'hc80;
    rom[2780 ] = 12'hc80;
    rom[2781 ] = 12'hc80;
    rom[2782 ] = 12'hc80;
    rom[2783 ] = 12'h000;
    rom[2784 ] = 12'h000;
    rom[2785 ] = 12'h000;
    rom[2786 ] = 12'h000;
    rom[2787 ] = 12'h000;
    rom[2788 ] = 12'h000;
    rom[2789 ] = 12'h000;
    rom[2790 ] = 12'h000;
    rom[2791 ] = 12'h000;
    rom[2792 ] = 12'h000;
    rom[2793 ] = 12'h000;
    rom[2794 ] = 12'h000;
    rom[2795 ] = 12'h000;
    rom[2796 ] = 12'h000;
    rom[2797 ] = 12'h000;
    rom[2798 ] = 12'h000;
    rom[2799 ] = 12'h000;
    rom[2800 ] = 12'h000;
    rom[2801 ] = 12'h000;
    rom[2802 ] = 12'h000;
    rom[2803 ] = 12'h000;
    rom[2804 ] = 12'h000;
    rom[2805 ] = 12'h000;
    rom[2806 ] = 12'h000;
    rom[2807 ] = 12'h000;
    rom[2808 ] = 12'h000;
    rom[2809 ] = 12'h000;
    rom[2810 ] = 12'h000;
    rom[2811 ] = 12'h000;
    rom[2812 ] = 12'h000;
    rom[2813 ] = 12'h000;
    rom[2814 ] = 12'h000;
    rom[2815 ] = 12'h000;
    rom[2816 ] = 12'h000;
    rom[2817 ] = 12'h000;
    rom[2818 ] = 12'h000;
    rom[2819 ] = 12'h000;
    rom[2820 ] = 12'h000;
    rom[2821 ] = 12'h000;
    rom[2822 ] = 12'h000;
    rom[2823 ] = 12'h000;
    rom[2824 ] = 12'h000;
    rom[2825 ] = 12'h000;
    rom[2826 ] = 12'h000;
    rom[2827 ] = 12'h000;
    rom[2828 ] = 12'h000;
    rom[2829 ] = 12'h000;
    rom[2830 ] = 12'h000;
    rom[2831 ] = 12'hea0;
    rom[2832 ] = 12'hea0;
    rom[2833 ] = 12'hea0;
    rom[2834 ] = 12'hea0;
    rom[2835 ] = 12'hea0;
    rom[2836 ] = 12'hea0;
    rom[2837 ] = 12'hea0;
    rom[2838 ] = 12'hea0;
    rom[2839 ] = 12'hea0;
    rom[2840 ] = 12'hea0;
    rom[2841 ] = 12'hea0;
    rom[2842 ] = 12'hea0;
    rom[2843 ] = 12'hea0;
    rom[2844 ] = 12'hea0;
    rom[2845 ] = 12'hea0;
    rom[2846 ] = 12'hea0;
    rom[2847 ] = 12'hea0;
    rom[2848 ] = 12'hea0;
    rom[2849 ] = 12'hea0;
    rom[2850 ] = 12'hea0;
    rom[2851 ] = 12'hea0;
    rom[2852 ] = 12'hea0;
    rom[2853 ] = 12'hea0;
    rom[2854 ] = 12'h000;
    rom[2855 ] = 12'h000;
    rom[2856 ] = 12'h000;
    rom[2857 ] = 12'h000;
    rom[2858 ] = 12'h000;
    rom[2859 ] = 12'h000;
    rom[2860 ] = 12'h000;
    rom[2861 ] = 12'h000;
    rom[2862 ] = 12'h000;
    rom[2863 ] = 12'h000;
    rom[2864 ] = 12'h000;
    rom[2865 ] = 12'h000;
    rom[2866 ] = 12'h000;
    rom[2867 ] = 12'h000;
    rom[2868 ] = 12'h000;
    rom[2869 ] = 12'h000;
    rom[2870 ] = 12'h000;
    rom[2871 ] = 12'h000;
    rom[2872 ] = 12'h000;
    rom[2873 ] = 12'h000;
    rom[2874 ] = 12'h000;
    rom[2875 ] = 12'h000;
    rom[2876 ] = 12'h000;
    rom[2877 ] = 12'h000;
    rom[2878 ] = 12'h000;
    rom[2879 ] = 12'h000;
    rom[2880 ] = 12'h000;
    rom[2881 ] = 12'h000;
    rom[2882 ] = 12'h000;
    rom[2883 ] = 12'h000;
    rom[2884 ] = 12'h000;
    rom[2885 ] = 12'h000;
    rom[2886 ] = 12'h000;
    rom[2887 ] = 12'h000;
    rom[2888 ] = 12'h000;
    rom[2889 ] = 12'h000;
    rom[2890 ] = 12'h000;
    rom[2891 ] = 12'h000;
    rom[2892 ] = 12'h000;
    rom[2893 ] = 12'h000;
    rom[2894 ] = 12'h000;
    rom[2895 ] = 12'h000;
    rom[2896 ] = 12'h000;
    rom[2897 ] = 12'h000;
    rom[2898 ] = 12'h000;
    rom[2899 ] = 12'h000;
    rom[2900 ] = 12'h000;
    rom[2901 ] = 12'h000;
    rom[2902 ] = 12'h000;
    rom[2903 ] = 12'h000;
    rom[2904 ] = 12'h000;
    rom[2905 ] = 12'h000;
    rom[2906 ] = 12'hc80;
    rom[2907 ] = 12'hc80;
    rom[2908 ] = 12'hc80;
    rom[2909 ] = 12'h000;
    rom[2910 ] = 12'h000;
    rom[2911 ] = 12'h000;
    rom[2912 ] = 12'h000;
    rom[2913 ] = 12'h000;
    rom[2914 ] = 12'h000;
    rom[2915 ] = 12'h000;
    rom[2916 ] = 12'h000;
    rom[2917 ] = 12'h000;
    rom[2918 ] = 12'h000;
    rom[2919 ] = 12'h000;
    rom[2920 ] = 12'h000;
    rom[2921 ] = 12'h000;
    rom[2922 ] = 12'h000;
    rom[2923 ] = 12'h000;
    rom[2924 ] = 12'h000;
    rom[2925 ] = 12'h000;
    rom[2926 ] = 12'h000;
    rom[2927 ] = 12'h000;
    rom[2928 ] = 12'h000;
    rom[2929 ] = 12'h000;
    rom[2930 ] = 12'h000;
    rom[2931 ] = 12'h000;
    rom[2932 ] = 12'h000;
    rom[2933 ] = 12'h000;
    rom[2934 ] = 12'h000;
    rom[2935 ] = 12'h000;
    rom[2936 ] = 12'h000;
    rom[2937 ] = 12'h000;
    rom[2938 ] = 12'h000;
    rom[2939 ] = 12'h000;
    rom[2940 ] = 12'h000;
    rom[2941 ] = 12'h000;
    rom[2942 ] = 12'h000;
    rom[2943 ] = 12'h000;
    rom[2944 ] = 12'h000;
    rom[2945 ] = 12'h000;
    rom[2946 ] = 12'h000;
    rom[2947 ] = 12'h000;
    rom[2948 ] = 12'h000;
    rom[2949 ] = 12'h000;
    rom[2950 ] = 12'h000;
    rom[2951 ] = 12'h000;
    rom[2952 ] = 12'h000;
    rom[2953 ] = 12'h000;
    rom[2954 ] = 12'h000;
    rom[2955 ] = 12'h000;
    rom[2956 ] = 12'h000;
    rom[2957 ] = 12'h000;
    rom[2958 ] = 12'hdb1;
    rom[2959 ] = 12'hda1;
    rom[2960 ] = 12'hda1;
    rom[2961 ] = 12'hea0;
    rom[2962 ] = 12'hea0;
    rom[2963 ] = 12'hea0;
    rom[2964 ] = 12'hea0;
    rom[2965 ] = 12'hea0;
    rom[2966 ] = 12'hea0;
    rom[2967 ] = 12'hea0;
    rom[2968 ] = 12'hea0;
    rom[2969 ] = 12'hea0;
    rom[2970 ] = 12'hea0;
    rom[2971 ] = 12'hea0;
    rom[2972 ] = 12'hea0;
    rom[2973 ] = 12'hea0;
    rom[2974 ] = 12'hea0;
    rom[2975 ] = 12'hea0;
    rom[2976 ] = 12'hea0;
    rom[2977 ] = 12'hea0;
    rom[2978 ] = 12'hea0;
    rom[2979 ] = 12'hea0;
    rom[2980 ] = 12'hfa0;
    rom[2981 ] = 12'h000;
    rom[2982 ] = 12'h000;
    rom[2983 ] = 12'h000;
    rom[2984 ] = 12'h000;
    rom[2985 ] = 12'h000;
    rom[2986 ] = 12'h000;
    rom[2987 ] = 12'h000;
    rom[2988 ] = 12'h000;
    rom[2989 ] = 12'h000;
    rom[2990 ] = 12'h000;
    rom[2991 ] = 12'h000;
    rom[2992 ] = 12'h000;
    rom[2993 ] = 12'h000;
    rom[2994 ] = 12'h000;
    rom[2995 ] = 12'h000;
    rom[2996 ] = 12'h000;
    rom[2997 ] = 12'h000;
    rom[2998 ] = 12'h000;
    rom[2999 ] = 12'h000;
    rom[3000 ] = 12'h000;
    rom[3001 ] = 12'h000;
    rom[3002 ] = 12'h000;
    rom[3003 ] = 12'h000;
    rom[3004 ] = 12'h000;
    rom[3005 ] = 12'h000;
    rom[3006 ] = 12'h000;
    rom[3007 ] = 12'h000;
    rom[3008 ] = 12'h000;
    rom[3009 ] = 12'h000;
    rom[3010 ] = 12'h000;
    rom[3011 ] = 12'h000;
    rom[3012 ] = 12'h000;
    rom[3013 ] = 12'h000;
    rom[3014 ] = 12'h000;
    rom[3015 ] = 12'h000;
    rom[3016 ] = 12'h000;
    rom[3017 ] = 12'h000;
    rom[3018 ] = 12'h000;
    rom[3019 ] = 12'h000;
    rom[3020 ] = 12'h000;
    rom[3021 ] = 12'h000;
    rom[3022 ] = 12'h000;
    rom[3023 ] = 12'h000;
    rom[3024 ] = 12'h000;
    rom[3025 ] = 12'h000;
    rom[3026 ] = 12'h000;
    rom[3027 ] = 12'h000;
    rom[3028 ] = 12'h000;
    rom[3029 ] = 12'h000;
    rom[3030 ] = 12'h000;
    rom[3031 ] = 12'h000;
    rom[3032 ] = 12'h000;
    rom[3033 ] = 12'h000;
    rom[3034 ] = 12'h000;
    rom[3035 ] = 12'hc80;
    rom[3036 ] = 12'h000;
    rom[3037 ] = 12'h000;
    rom[3038 ] = 12'h000;
    rom[3039 ] = 12'h000;
    rom[3040 ] = 12'h000;
    rom[3041 ] = 12'h000;
    rom[3042 ] = 12'h000;
    rom[3043 ] = 12'h000;
    rom[3044 ] = 12'h000;
    rom[3045 ] = 12'h000;
    rom[3046 ] = 12'h000;
    rom[3047 ] = 12'h000;
    rom[3048 ] = 12'h000;
    rom[3049 ] = 12'h000;
    rom[3050 ] = 12'h000;
    rom[3051 ] = 12'h000;
    rom[3052 ] = 12'h000;
    rom[3053 ] = 12'h000;
    rom[3054 ] = 12'h000;
    rom[3055 ] = 12'h000;
    rom[3056 ] = 12'h000;
    rom[3057 ] = 12'h000;
    rom[3058 ] = 12'h000;
    rom[3059 ] = 12'h000;
    rom[3060 ] = 12'h000;
    rom[3061 ] = 12'h000;
    rom[3062 ] = 12'h000;
    rom[3063 ] = 12'h000;
    rom[3064 ] = 12'h000;
    rom[3065 ] = 12'h000;
    rom[3066 ] = 12'h000;
    rom[3067 ] = 12'h000;
    rom[3068 ] = 12'h000;
    rom[3069 ] = 12'h000;
    rom[3070 ] = 12'h000;
    rom[3071 ] = 12'h000;
    rom[3072 ] = 12'h000;
    rom[3073 ] = 12'h000;
    rom[3074 ] = 12'h000;
    rom[3075 ] = 12'h000;
    rom[3076 ] = 12'h000;
    rom[3077 ] = 12'h000;
    rom[3078 ] = 12'h000;
    rom[3079 ] = 12'h000;
    rom[3080 ] = 12'h000;
    rom[3081 ] = 12'h000;
    rom[3082 ] = 12'h000;
    rom[3083 ] = 12'h000;
    rom[3084 ] = 12'h000;
    rom[3085 ] = 12'h000;
    rom[3086 ] = 12'hda1;
    rom[3087 ] = 12'hda1;
    rom[3088 ] = 12'hda1;
    rom[3089 ] = 12'hda1;
    rom[3090 ] = 12'hda1;
    rom[3091 ] = 12'hda1;
    rom[3092 ] = 12'hea0;
    rom[3093 ] = 12'hea0;
    rom[3094 ] = 12'hea0;
    rom[3095 ] = 12'hea0;
    rom[3096 ] = 12'hea0;
    rom[3097 ] = 12'hea0;
    rom[3098 ] = 12'hea0;
    rom[3099 ] = 12'hea0;
    rom[3100 ] = 12'hea0;
    rom[3101 ] = 12'hea0;
    rom[3102 ] = 12'hea0;
    rom[3103 ] = 12'hea0;
    rom[3104 ] = 12'hea0;
    rom[3105 ] = 12'hea0;
    rom[3106 ] = 12'hea0;
    rom[3107 ] = 12'h000;
    rom[3108 ] = 12'h000;
    rom[3109 ] = 12'h000;
    rom[3110 ] = 12'h000;
    rom[3111 ] = 12'h000;
    rom[3112 ] = 12'h000;
    rom[3113 ] = 12'h000;
    rom[3114 ] = 12'h000;
    rom[3115 ] = 12'h000;
    rom[3116 ] = 12'h000;
    rom[3117 ] = 12'h000;
    rom[3118 ] = 12'h000;
    rom[3119 ] = 12'h000;
    rom[3120 ] = 12'h000;
    rom[3121 ] = 12'h000;
    rom[3122 ] = 12'h000;
    rom[3123 ] = 12'h000;
    rom[3124 ] = 12'h000;
    rom[3125 ] = 12'h000;
    rom[3126 ] = 12'h000;
    rom[3127 ] = 12'h000;
    rom[3128 ] = 12'h000;
    rom[3129 ] = 12'h000;
    rom[3130 ] = 12'h000;
    rom[3131 ] = 12'h000;
    rom[3132 ] = 12'h000;
    rom[3133 ] = 12'h000;
    rom[3134 ] = 12'h000;
    rom[3135 ] = 12'h000;
    rom[3136 ] = 12'h000;
    rom[3137 ] = 12'h000;
    rom[3138 ] = 12'h000;
    rom[3139 ] = 12'h000;
    rom[3140 ] = 12'h000;
    rom[3141 ] = 12'h000;
    rom[3142 ] = 12'h000;
    rom[3143 ] = 12'h000;
    rom[3144 ] = 12'h000;
    rom[3145 ] = 12'h000;
    rom[3146 ] = 12'h000;
    rom[3147 ] = 12'h000;
    rom[3148 ] = 12'h000;
    rom[3149 ] = 12'h000;
    rom[3150 ] = 12'h000;
    rom[3151 ] = 12'h000;
    rom[3152 ] = 12'h000;
    rom[3153 ] = 12'h000;
    rom[3154 ] = 12'h000;
    rom[3155 ] = 12'h000;
    rom[3156 ] = 12'h000;
    rom[3157 ] = 12'h000;
    rom[3158 ] = 12'h000;
    rom[3159 ] = 12'h000;
    rom[3160 ] = 12'h000;
    rom[3161 ] = 12'h000;
    rom[3162 ] = 12'h000;
    rom[3163 ] = 12'h000;
    rom[3164 ] = 12'h000;
    rom[3165 ] = 12'h000;
    rom[3166 ] = 12'h000;
    rom[3167 ] = 12'h000;
    rom[3168 ] = 12'h000;
    rom[3169 ] = 12'h000;
    rom[3170 ] = 12'h000;
    rom[3171 ] = 12'h000;
    rom[3172 ] = 12'h000;
    rom[3173 ] = 12'h000;
    rom[3174 ] = 12'h000;
    rom[3175 ] = 12'h000;
    rom[3176 ] = 12'h000;
    rom[3177 ] = 12'h000;
    rom[3178 ] = 12'h000;
    rom[3179 ] = 12'h000;
    rom[3180 ] = 12'h000;
    rom[3181 ] = 12'h000;
    rom[3182 ] = 12'h000;
    rom[3183 ] = 12'h000;
    rom[3184 ] = 12'h000;
    rom[3185 ] = 12'h000;
    rom[3186 ] = 12'h000;
    rom[3187 ] = 12'h000;
    rom[3188 ] = 12'h000;
    rom[3189 ] = 12'h000;
    rom[3190 ] = 12'h000;
    rom[3191 ] = 12'h000;
    rom[3192 ] = 12'h000;
    rom[3193 ] = 12'h000;
    rom[3194 ] = 12'h000;
    rom[3195 ] = 12'h000;
    rom[3196 ] = 12'h000;
    rom[3197 ] = 12'h000;
    rom[3198 ] = 12'h000;
    rom[3199 ] = 12'h000;
    rom[3200 ] = 12'h000;
    rom[3201 ] = 12'h000;
    rom[3202 ] = 12'h000;
    rom[3203 ] = 12'h000;
    rom[3204 ] = 12'h000;
    rom[3205 ] = 12'h000;
    rom[3206 ] = 12'h000;
    rom[3207 ] = 12'h000;
    rom[3208 ] = 12'h000;
    rom[3209 ] = 12'h000;
    rom[3210 ] = 12'h000;
    rom[3211 ] = 12'h000;
    rom[3212 ] = 12'h000;
    rom[3213 ] = 12'hda1;
    rom[3214 ] = 12'hda1;
    rom[3215 ] = 12'hda1;
    rom[3216 ] = 12'hda1;
    rom[3217 ] = 12'hda1;
    rom[3218 ] = 12'hda1;
    rom[3219 ] = 12'hda1;
    rom[3220 ] = 12'hda1;
    rom[3221 ] = 12'hda1;
    rom[3222 ] = 12'hea0;
    rom[3223 ] = 12'hea0;
    rom[3224 ] = 12'hea0;
    rom[3225 ] = 12'hea0;
    rom[3226 ] = 12'hea0;
    rom[3227 ] = 12'hea0;
    rom[3228 ] = 12'hea0;
    rom[3229 ] = 12'hea0;
    rom[3230 ] = 12'hea0;
    rom[3231 ] = 12'hea0;
    rom[3232 ] = 12'hea0;
    rom[3233 ] = 12'hea0;
    rom[3234 ] = 12'h000;
    rom[3235 ] = 12'h000;
    rom[3236 ] = 12'h000;
    rom[3237 ] = 12'h000;
    rom[3238 ] = 12'h000;
    rom[3239 ] = 12'h000;
    rom[3240 ] = 12'h000;
    rom[3241 ] = 12'h000;
    rom[3242 ] = 12'h000;
    rom[3243 ] = 12'h000;
    rom[3244 ] = 12'h000;
    rom[3245 ] = 12'h000;
    rom[3246 ] = 12'h000;
    rom[3247 ] = 12'h000;
    rom[3248 ] = 12'h000;
    rom[3249 ] = 12'h000;
    rom[3250 ] = 12'h000;
    rom[3251 ] = 12'h000;
    rom[3252 ] = 12'h000;
    rom[3253 ] = 12'h000;
    rom[3254 ] = 12'h000;
    rom[3255 ] = 12'h000;
    rom[3256 ] = 12'h000;
    rom[3257 ] = 12'h000;
    rom[3258 ] = 12'h000;
    rom[3259 ] = 12'h000;
    rom[3260 ] = 12'h000;
    rom[3261 ] = 12'h000;
    rom[3262 ] = 12'h000;
    rom[3263 ] = 12'h000;
    rom[3264 ] = 12'h000;
    rom[3265 ] = 12'h000;
    rom[3266 ] = 12'h000;
    rom[3267 ] = 12'h000;
    rom[3268 ] = 12'h000;
    rom[3269 ] = 12'h000;
    rom[3270 ] = 12'h000;
    rom[3271 ] = 12'h000;
    rom[3272 ] = 12'h000;
    rom[3273 ] = 12'h000;
    rom[3274 ] = 12'h000;
    rom[3275 ] = 12'h000;
    rom[3276 ] = 12'h000;
    rom[3277 ] = 12'h000;
    rom[3278 ] = 12'h000;
    rom[3279 ] = 12'h000;
    rom[3280 ] = 12'h000;
    rom[3281 ] = 12'h000;
    rom[3282 ] = 12'h000;
    rom[3283 ] = 12'h000;
    rom[3284 ] = 12'h000;
    rom[3285 ] = 12'h000;
    rom[3286 ] = 12'h000;
    rom[3287 ] = 12'h000;
    rom[3288 ] = 12'h000;
    rom[3289 ] = 12'h000;
    rom[3290 ] = 12'h000;
    rom[3291 ] = 12'h000;
    rom[3292 ] = 12'h000;
    rom[3293 ] = 12'h000;
    rom[3294 ] = 12'h000;
    rom[3295 ] = 12'h000;
    rom[3296 ] = 12'h000;
    rom[3297 ] = 12'h000;
    rom[3298 ] = 12'h000;
    rom[3299 ] = 12'h000;
    rom[3300 ] = 12'h000;
    rom[3301 ] = 12'h000;
    rom[3302 ] = 12'h000;
    rom[3303 ] = 12'h000;
    rom[3304 ] = 12'h000;
    rom[3305 ] = 12'h000;
    rom[3306 ] = 12'h000;
    rom[3307 ] = 12'h000;
    rom[3308 ] = 12'h000;
    rom[3309 ] = 12'h000;
    rom[3310 ] = 12'h000;
    rom[3311 ] = 12'h000;
    rom[3312 ] = 12'h000;
    rom[3313 ] = 12'h000;
    rom[3314 ] = 12'h3a2;
    rom[3315 ] = 12'h000;
    rom[3316 ] = 12'h000;
    rom[3317 ] = 12'h000;
    rom[3318 ] = 12'h000;
    rom[3319 ] = 12'h000;
    rom[3320 ] = 12'h000;
    rom[3321 ] = 12'h000;
    rom[3322 ] = 12'h000;
    rom[3323 ] = 12'h000;
    rom[3324 ] = 12'h000;
    rom[3325 ] = 12'h000;
    rom[3326 ] = 12'h000;
    rom[3327 ] = 12'h000;
    rom[3328 ] = 12'h000;
    rom[3329 ] = 12'h000;
    rom[3330 ] = 12'h000;
    rom[3331 ] = 12'h000;
    rom[3332 ] = 12'h000;
    rom[3333 ] = 12'h000;
    rom[3334 ] = 12'h000;
    rom[3335 ] = 12'h000;
    rom[3336 ] = 12'h000;
    rom[3337 ] = 12'h000;
    rom[3338 ] = 12'h000;
    rom[3339 ] = 12'h000;
    rom[3340 ] = 12'hca2;
    rom[3341 ] = 12'hca1;
    rom[3342 ] = 12'hca1;
    rom[3343 ] = 12'hda1;
    rom[3344 ] = 12'hda1;
    rom[3345 ] = 12'hda1;
    rom[3346 ] = 12'hda1;
    rom[3347 ] = 12'hda1;
    rom[3348 ] = 12'hda1;
    rom[3349 ] = 12'hda1;
    rom[3350 ] = 12'hda1;
    rom[3351 ] = 12'hda1;
    rom[3352 ] = 12'hda1;
    rom[3353 ] = 12'hea0;
    rom[3354 ] = 12'hea0;
    rom[3355 ] = 12'hea0;
    rom[3356 ] = 12'hea0;
    rom[3357 ] = 12'hea0;
    rom[3358 ] = 12'hea0;
    rom[3359 ] = 12'hea0;
    rom[3360 ] = 12'hea0;
    rom[3361 ] = 12'h000;
    rom[3362 ] = 12'h000;
    rom[3363 ] = 12'h000;
    rom[3364 ] = 12'h000;
    rom[3365 ] = 12'h000;
    rom[3366 ] = 12'h000;
    rom[3367 ] = 12'h000;
    rom[3368 ] = 12'h000;
    rom[3369 ] = 12'h000;
    rom[3370 ] = 12'h000;
    rom[3371 ] = 12'h000;
    rom[3372 ] = 12'h000;
    rom[3373 ] = 12'h000;
    rom[3374 ] = 12'h000;
    rom[3375 ] = 12'h000;
    rom[3376 ] = 12'h000;
    rom[3377 ] = 12'h000;
    rom[3378 ] = 12'h000;
    rom[3379 ] = 12'h000;
    rom[3380 ] = 12'h000;
    rom[3381 ] = 12'h000;
    rom[3382 ] = 12'h000;
    rom[3383 ] = 12'h000;
    rom[3384 ] = 12'h000;
    rom[3385 ] = 12'h000;
    rom[3386 ] = 12'h000;
    rom[3387 ] = 12'h000;
    rom[3388 ] = 12'h000;
    rom[3389 ] = 12'h000;
    rom[3390 ] = 12'h000;
    rom[3391 ] = 12'h000;
    rom[3392 ] = 12'h000;
    rom[3393 ] = 12'h000;
    rom[3394 ] = 12'h000;
    rom[3395 ] = 12'h000;
    rom[3396 ] = 12'h000;
    rom[3397 ] = 12'h000;
    rom[3398 ] = 12'h000;
    rom[3399 ] = 12'h000;
    rom[3400 ] = 12'h000;
    rom[3401 ] = 12'h000;
    rom[3402 ] = 12'h000;
    rom[3403 ] = 12'h000;
    rom[3404 ] = 12'h000;
    rom[3405 ] = 12'h000;
    rom[3406 ] = 12'h000;
    rom[3407 ] = 12'h000;
    rom[3408 ] = 12'h000;
    rom[3409 ] = 12'h000;
    rom[3410 ] = 12'h000;
    rom[3411 ] = 12'h000;
    rom[3412 ] = 12'h000;
    rom[3413 ] = 12'h000;
    rom[3414 ] = 12'h000;
    rom[3415 ] = 12'h000;
    rom[3416 ] = 12'h000;
    rom[3417 ] = 12'h000;
    rom[3418 ] = 12'h000;
    rom[3419 ] = 12'h000;
    rom[3420 ] = 12'h000;
    rom[3421 ] = 12'h000;
    rom[3422 ] = 12'h000;
    rom[3423 ] = 12'h000;
    rom[3424 ] = 12'h000;
    rom[3425 ] = 12'h000;
    rom[3426 ] = 12'h000;
    rom[3427 ] = 12'h000;
    rom[3428 ] = 12'h000;
    rom[3429 ] = 12'h000;
    rom[3430 ] = 12'h000;
    rom[3431 ] = 12'h000;
    rom[3432 ] = 12'h000;
    rom[3433 ] = 12'h000;
    rom[3434 ] = 12'h000;
    rom[3435 ] = 12'h000;
    rom[3436 ] = 12'h000;
    rom[3437 ] = 12'h000;
    rom[3438 ] = 12'h000;
    rom[3439 ] = 12'h000;
    rom[3440 ] = 12'h3a1;
    rom[3441 ] = 12'h3a2;
    rom[3442 ] = 12'h3a2;
    rom[3443 ] = 12'h3a2;
    rom[3444 ] = 12'h000;
    rom[3445 ] = 12'h000;
    rom[3446 ] = 12'h000;
    rom[3447 ] = 12'h000;
    rom[3448 ] = 12'h000;
    rom[3449 ] = 12'h000;
    rom[3450 ] = 12'h000;
    rom[3451 ] = 12'h000;
    rom[3452 ] = 12'h000;
    rom[3453 ] = 12'h000;
    rom[3454 ] = 12'h000;
    rom[3455 ] = 12'h000;
    rom[3456 ] = 12'h000;
    rom[3457 ] = 12'h000;
    rom[3458 ] = 12'h000;
    rom[3459 ] = 12'h000;
    rom[3460 ] = 12'h000;
    rom[3461 ] = 12'h000;
    rom[3462 ] = 12'h000;
    rom[3463 ] = 12'h000;
    rom[3464 ] = 12'h000;
    rom[3465 ] = 12'h000;
    rom[3466 ] = 12'h000;
    rom[3467 ] = 12'hca2;
    rom[3468 ] = 12'hca2;
    rom[3469 ] = 12'hca2;
    rom[3470 ] = 12'hca2;
    rom[3471 ] = 12'hca2;
    rom[3472 ] = 12'hca1;
    rom[3473 ] = 12'hda1;
    rom[3474 ] = 12'hda1;
    rom[3475 ] = 12'hda1;
    rom[3476 ] = 12'hda1;
    rom[3477 ] = 12'hda1;
    rom[3478 ] = 12'hda1;
    rom[3479 ] = 12'hda1;
    rom[3480 ] = 12'hda1;
    rom[3481 ] = 12'hda1;
    rom[3482 ] = 12'hda1;
    rom[3483 ] = 12'hea0;
    rom[3484 ] = 12'hea0;
    rom[3485 ] = 12'hea0;
    rom[3486 ] = 12'hea0;
    rom[3487 ] = 12'h000;
    rom[3488 ] = 12'h000;
    rom[3489 ] = 12'h000;
    rom[3490 ] = 12'h000;
    rom[3491 ] = 12'h000;
    rom[3492 ] = 12'h000;
    rom[3493 ] = 12'h000;
    rom[3494 ] = 12'h000;
    rom[3495 ] = 12'h000;
    rom[3496 ] = 12'h000;
    rom[3497 ] = 12'h000;
    rom[3498 ] = 12'h000;
    rom[3499 ] = 12'h000;
    rom[3500 ] = 12'h000;
    rom[3501 ] = 12'h000;
    rom[3502 ] = 12'h000;
    rom[3503 ] = 12'h000;
    rom[3504 ] = 12'h000;
    rom[3505 ] = 12'h000;
    rom[3506 ] = 12'h000;
    rom[3507 ] = 12'h000;
    rom[3508 ] = 12'h000;
    rom[3509 ] = 12'h000;
    rom[3510 ] = 12'h000;
    rom[3511 ] = 12'h000;
    rom[3512 ] = 12'h000;
    rom[3513 ] = 12'h000;
    rom[3514 ] = 12'h000;
    rom[3515 ] = 12'h000;
    rom[3516 ] = 12'h000;
    rom[3517 ] = 12'h000;
    rom[3518 ] = 12'h000;
    rom[3519 ] = 12'h000;
    rom[3520 ] = 12'h000;
    rom[3521 ] = 12'h000;
    rom[3522 ] = 12'h000;
    rom[3523 ] = 12'h000;
    rom[3524 ] = 12'h000;
    rom[3525 ] = 12'h000;
    rom[3526 ] = 12'h000;
    rom[3527 ] = 12'h000;
    rom[3528 ] = 12'h000;
    rom[3529 ] = 12'h000;
    rom[3530 ] = 12'h000;
    rom[3531 ] = 12'h000;
    rom[3532 ] = 12'h000;
    rom[3533 ] = 12'h000;
    rom[3534 ] = 12'h000;
    rom[3535 ] = 12'h000;
    rom[3536 ] = 12'h000;
    rom[3537 ] = 12'h000;
    rom[3538 ] = 12'h000;
    rom[3539 ] = 12'h000;
    rom[3540 ] = 12'h000;
    rom[3541 ] = 12'h000;
    rom[3542 ] = 12'h000;
    rom[3543 ] = 12'h000;
    rom[3544 ] = 12'h000;
    rom[3545 ] = 12'h000;
    rom[3546 ] = 12'h000;
    rom[3547 ] = 12'h000;
    rom[3548 ] = 12'h000;
    rom[3549 ] = 12'h000;
    rom[3550 ] = 12'h000;
    rom[3551 ] = 12'h000;
    rom[3552 ] = 12'h000;
    rom[3553 ] = 12'h000;
    rom[3554 ] = 12'h000;
    rom[3555 ] = 12'h000;
    rom[3556 ] = 12'h000;
    rom[3557 ] = 12'h000;
    rom[3558 ] = 12'h000;
    rom[3559 ] = 12'h000;
    rom[3560 ] = 12'h000;
    rom[3561 ] = 12'h000;
    rom[3562 ] = 12'h000;
    rom[3563 ] = 12'h000;
    rom[3564 ] = 12'h000;
    rom[3565 ] = 12'h000;
    rom[3566 ] = 12'h000;
    rom[3567 ] = 12'h3a2;
    rom[3568 ] = 12'h3a2;
    rom[3569 ] = 12'h3a2;
    rom[3570 ] = 12'h3a2;
    rom[3571 ] = 12'h3a2;
    rom[3572 ] = 12'h392;
    rom[3573 ] = 12'h000;
    rom[3574 ] = 12'h000;
    rom[3575 ] = 12'h000;
    rom[3576 ] = 12'h000;
    rom[3577 ] = 12'h000;
    rom[3578 ] = 12'h000;
    rom[3579 ] = 12'h000;
    rom[3580 ] = 12'h000;
    rom[3581 ] = 12'h000;
    rom[3582 ] = 12'h000;
    rom[3583 ] = 12'h000;
    rom[3584 ] = 12'h000;
    rom[3585 ] = 12'h000;
    rom[3586 ] = 12'h000;
    rom[3587 ] = 12'h000;
    rom[3588 ] = 12'h000;
    rom[3589 ] = 12'h000;
    rom[3590 ] = 12'h000;
    rom[3591 ] = 12'h000;
    rom[3592 ] = 12'h000;
    rom[3593 ] = 12'h000;
    rom[3594 ] = 12'h000;
    rom[3595 ] = 12'hca2;
    rom[3596 ] = 12'hca2;
    rom[3597 ] = 12'hca2;
    rom[3598 ] = 12'hca2;
    rom[3599 ] = 12'hca2;
    rom[3600 ] = 12'hca2;
    rom[3601 ] = 12'hca2;
    rom[3602 ] = 12'hca1;
    rom[3603 ] = 12'hca1;
    rom[3604 ] = 12'hda1;
    rom[3605 ] = 12'hda1;
    rom[3606 ] = 12'hda1;
    rom[3607 ] = 12'hda1;
    rom[3608 ] = 12'hda1;
    rom[3609 ] = 12'hda1;
    rom[3610 ] = 12'hda1;
    rom[3611 ] = 12'hda1;
    rom[3612 ] = 12'hda1;
    rom[3613 ] = 12'hda1;
    rom[3614 ] = 12'h000;
    rom[3615 ] = 12'h000;
    rom[3616 ] = 12'h000;
    rom[3617 ] = 12'h000;
    rom[3618 ] = 12'h000;
    rom[3619 ] = 12'h000;
    rom[3620 ] = 12'h000;
    rom[3621 ] = 12'h000;
    rom[3622 ] = 12'h000;
    rom[3623 ] = 12'h000;
    rom[3624 ] = 12'h000;
    rom[3625 ] = 12'h000;
    rom[3626 ] = 12'h000;
    rom[3627 ] = 12'h000;
    rom[3628 ] = 12'h000;
    rom[3629 ] = 12'h000;
    rom[3630 ] = 12'h000;
    rom[3631 ] = 12'h000;
    rom[3632 ] = 12'h000;
    rom[3633 ] = 12'h000;
    rom[3634 ] = 12'h000;
    rom[3635 ] = 12'h000;
    rom[3636 ] = 12'h000;
    rom[3637 ] = 12'h000;
    rom[3638 ] = 12'h000;
    rom[3639 ] = 12'h000;
    rom[3640 ] = 12'h000;
    rom[3641 ] = 12'h000;
    rom[3642 ] = 12'h000;
    rom[3643 ] = 12'h000;
    rom[3644 ] = 12'h000;
    rom[3645 ] = 12'h000;
    rom[3646 ] = 12'h000;
    rom[3647 ] = 12'h000;
    rom[3648 ] = 12'h000;
    rom[3649 ] = 12'h000;
    rom[3650 ] = 12'h000;
    rom[3651 ] = 12'h000;
    rom[3652 ] = 12'h000;
    rom[3653 ] = 12'h000;
    rom[3654 ] = 12'h000;
    rom[3655 ] = 12'h000;
    rom[3656 ] = 12'h000;
    rom[3657 ] = 12'h000;
    rom[3658 ] = 12'h000;
    rom[3659 ] = 12'h000;
    rom[3660 ] = 12'h000;
    rom[3661 ] = 12'h000;
    rom[3662 ] = 12'h000;
    rom[3663 ] = 12'h000;
    rom[3664 ] = 12'h000;
    rom[3665 ] = 12'h000;
    rom[3666 ] = 12'h000;
    rom[3667 ] = 12'h000;
    rom[3668 ] = 12'h000;
    rom[3669 ] = 12'h000;
    rom[3670 ] = 12'h000;
    rom[3671 ] = 12'h000;
    rom[3672 ] = 12'h000;
    rom[3673 ] = 12'h000;
    rom[3674 ] = 12'h000;
    rom[3675 ] = 12'h000;
    rom[3676 ] = 12'h000;
    rom[3677 ] = 12'h000;
    rom[3678 ] = 12'h000;
    rom[3679 ] = 12'h000;
    rom[3680 ] = 12'h000;
    rom[3681 ] = 12'h000;
    rom[3682 ] = 12'h000;
    rom[3683 ] = 12'h000;
    rom[3684 ] = 12'h000;
    rom[3685 ] = 12'h000;
    rom[3686 ] = 12'h000;
    rom[3687 ] = 12'h000;
    rom[3688 ] = 12'h000;
    rom[3689 ] = 12'h000;
    rom[3690 ] = 12'h000;
    rom[3691 ] = 12'h000;
    rom[3692 ] = 12'h000;
    rom[3693 ] = 12'h000;
    rom[3694 ] = 12'h3a2;
    rom[3695 ] = 12'h3a2;
    rom[3696 ] = 12'h3a2;
    rom[3697 ] = 12'h3a2;
    rom[3698 ] = 12'h3a2;
    rom[3699 ] = 12'h3a2;
    rom[3700 ] = 12'h3a2;
    rom[3701 ] = 12'h000;
    rom[3702 ] = 12'h000;
    rom[3703 ] = 12'h000;
    rom[3704 ] = 12'h000;
    rom[3705 ] = 12'h000;
    rom[3706 ] = 12'h000;
    rom[3707 ] = 12'h000;
    rom[3708 ] = 12'h000;
    rom[3709 ] = 12'h000;
    rom[3710 ] = 12'h000;
    rom[3711 ] = 12'h000;
    rom[3712 ] = 12'h000;
    rom[3713 ] = 12'h000;
    rom[3714 ] = 12'h000;
    rom[3715 ] = 12'h000;
    rom[3716 ] = 12'h000;
    rom[3717 ] = 12'h000;
    rom[3718 ] = 12'h000;
    rom[3719 ] = 12'h000;
    rom[3720 ] = 12'h000;
    rom[3721 ] = 12'h000;
    rom[3722 ] = 12'hbb2;
    rom[3723 ] = 12'hba2;
    rom[3724 ] = 12'hca2;
    rom[3725 ] = 12'hca2;
    rom[3726 ] = 12'hca2;
    rom[3727 ] = 12'hca2;
    rom[3728 ] = 12'hca2;
    rom[3729 ] = 12'hca2;
    rom[3730 ] = 12'hca2;
    rom[3731 ] = 12'hca2;
    rom[3732 ] = 12'hca2;
    rom[3733 ] = 12'hca1;
    rom[3734 ] = 12'hda1;
    rom[3735 ] = 12'hda1;
    rom[3736 ] = 12'hda1;
    rom[3737 ] = 12'hda1;
    rom[3738 ] = 12'hda1;
    rom[3739 ] = 12'hda1;
    rom[3740 ] = 12'hda1;
    rom[3741 ] = 12'h000;
    rom[3742 ] = 12'h000;
    rom[3743 ] = 12'h000;
    rom[3744 ] = 12'h000;
    rom[3745 ] = 12'h000;
    rom[3746 ] = 12'h000;
    rom[3747 ] = 12'h000;
    rom[3748 ] = 12'h000;
    rom[3749 ] = 12'h000;
    rom[3750 ] = 12'h000;
    rom[3751 ] = 12'h000;
    rom[3752 ] = 12'h000;
    rom[3753 ] = 12'h000;
    rom[3754 ] = 12'h000;
    rom[3755 ] = 12'h000;
    rom[3756 ] = 12'h000;
    rom[3757 ] = 12'h000;
    rom[3758 ] = 12'h000;
    rom[3759 ] = 12'h000;
    rom[3760 ] = 12'h000;
    rom[3761 ] = 12'h000;
    rom[3762 ] = 12'h000;
    rom[3763 ] = 12'h000;
    rom[3764 ] = 12'h000;
    rom[3765 ] = 12'h000;
    rom[3766 ] = 12'h000;
    rom[3767 ] = 12'h000;
    rom[3768 ] = 12'h000;
    rom[3769 ] = 12'h000;
    rom[3770 ] = 12'h000;
    rom[3771 ] = 12'h000;
    rom[3772 ] = 12'h000;
    rom[3773 ] = 12'h000;
    rom[3774 ] = 12'h000;
    rom[3775 ] = 12'h000;
    rom[3776 ] = 12'h000;
    rom[3777 ] = 12'h000;
    rom[3778 ] = 12'h000;
    rom[3779 ] = 12'h000;
    rom[3780 ] = 12'h000;
    rom[3781 ] = 12'h000;
    rom[3782 ] = 12'h000;
    rom[3783 ] = 12'h000;
    rom[3784 ] = 12'h000;
    rom[3785 ] = 12'h000;
    rom[3786 ] = 12'h000;
    rom[3787 ] = 12'h000;
    rom[3788 ] = 12'h000;
    rom[3789 ] = 12'h000;
    rom[3790 ] = 12'h000;
    rom[3791 ] = 12'h000;
    rom[3792 ] = 12'h000;
    rom[3793 ] = 12'h000;
    rom[3794 ] = 12'h000;
    rom[3795 ] = 12'h000;
    rom[3796 ] = 12'h000;
    rom[3797 ] = 12'h000;
    rom[3798 ] = 12'h000;
    rom[3799 ] = 12'h000;
    rom[3800 ] = 12'h000;
    rom[3801 ] = 12'h000;
    rom[3802 ] = 12'h000;
    rom[3803 ] = 12'h000;
    rom[3804 ] = 12'h000;
    rom[3805 ] = 12'h000;
    rom[3806 ] = 12'h000;
    rom[3807 ] = 12'h000;
    rom[3808 ] = 12'h000;
    rom[3809 ] = 12'h000;
    rom[3810 ] = 12'h000;
    rom[3811 ] = 12'h000;
    rom[3812 ] = 12'h000;
    rom[3813 ] = 12'h000;
    rom[3814 ] = 12'h000;
    rom[3815 ] = 12'h000;
    rom[3816 ] = 12'h000;
    rom[3817 ] = 12'h000;
    rom[3818 ] = 12'h000;
    rom[3819 ] = 12'h000;
    rom[3820 ] = 12'h3a2;
    rom[3821 ] = 12'h3a2;
    rom[3822 ] = 12'h3a2;
    rom[3823 ] = 12'h3a2;
    rom[3824 ] = 12'h3a2;
    rom[3825 ] = 12'h3a2;
    rom[3826 ] = 12'h3a2;
    rom[3827 ] = 12'h3a2;
    rom[3828 ] = 12'h3a2;
    rom[3829 ] = 12'h3a2;
    rom[3830 ] = 12'h000;
    rom[3831 ] = 12'h000;
    rom[3832 ] = 12'h000;
    rom[3833 ] = 12'h000;
    rom[3834 ] = 12'h000;
    rom[3835 ] = 12'h000;
    rom[3836 ] = 12'h000;
    rom[3837 ] = 12'h000;
    rom[3838 ] = 12'h000;
    rom[3839 ] = 12'h000;
    rom[3840 ] = 12'h000;
    rom[3841 ] = 12'h000;
    rom[3842 ] = 12'h000;
    rom[3843 ] = 12'h000;
    rom[3844 ] = 12'h000;
    rom[3845 ] = 12'h000;
    rom[3846 ] = 12'h000;
    rom[3847 ] = 12'h000;
    rom[3848 ] = 12'h000;
    rom[3849 ] = 12'hbb3;
    rom[3850 ] = 12'hbb3;
    rom[3851 ] = 12'hbb3;
    rom[3852 ] = 12'hbb2;
    rom[3853 ] = 12'hbb2;
    rom[3854 ] = 12'hba2;
    rom[3855 ] = 12'hca2;
    rom[3856 ] = 12'hca2;
    rom[3857 ] = 12'hca2;
    rom[3858 ] = 12'hca2;
    rom[3859 ] = 12'hca2;
    rom[3860 ] = 12'hca2;
    rom[3861 ] = 12'hca2;
    rom[3862 ] = 12'hca2;
    rom[3863 ] = 12'hca2;
    rom[3864 ] = 12'hca1;
    rom[3865 ] = 12'hda1;
    rom[3866 ] = 12'hda1;
    rom[3867 ] = 12'hda1;
    rom[3868 ] = 12'h000;
    rom[3869 ] = 12'h000;
    rom[3870 ] = 12'h000;
    rom[3871 ] = 12'h000;
    rom[3872 ] = 12'h000;
    rom[3873 ] = 12'h000;
    rom[3874 ] = 12'h000;
    rom[3875 ] = 12'h000;
    rom[3876 ] = 12'h000;
    rom[3877 ] = 12'h000;
    rom[3878 ] = 12'h000;
    rom[3879 ] = 12'h000;
    rom[3880 ] = 12'h000;
    rom[3881 ] = 12'h000;
    rom[3882 ] = 12'h000;
    rom[3883 ] = 12'h000;
    rom[3884 ] = 12'h000;
    rom[3885 ] = 12'h000;
    rom[3886 ] = 12'h000;
    rom[3887 ] = 12'h000;
    rom[3888 ] = 12'h000;
    rom[3889 ] = 12'h000;
    rom[3890 ] = 12'h000;
    rom[3891 ] = 12'h000;
    rom[3892 ] = 12'h000;
    rom[3893 ] = 12'h000;
    rom[3894 ] = 12'h000;
    rom[3895 ] = 12'h000;
    rom[3896 ] = 12'h000;
    rom[3897 ] = 12'h000;
    rom[3898 ] = 12'h000;
    rom[3899 ] = 12'h000;
    rom[3900 ] = 12'h000;
    rom[3901 ] = 12'h000;
    rom[3902 ] = 12'h000;
    rom[3903 ] = 12'h000;
    rom[3904 ] = 12'h000;
    rom[3905 ] = 12'h000;
    rom[3906 ] = 12'h000;
    rom[3907 ] = 12'h000;
    rom[3908 ] = 12'h000;
    rom[3909 ] = 12'h000;
    rom[3910 ] = 12'h000;
    rom[3911 ] = 12'h000;
    rom[3912 ] = 12'h000;
    rom[3913 ] = 12'h000;
    rom[3914 ] = 12'h000;
    rom[3915 ] = 12'h000;
    rom[3916 ] = 12'h000;
    rom[3917 ] = 12'h000;
    rom[3918 ] = 12'h000;
    rom[3919 ] = 12'h000;
    rom[3920 ] = 12'h000;
    rom[3921 ] = 12'h000;
    rom[3922 ] = 12'h000;
    rom[3923 ] = 12'h000;
    rom[3924 ] = 12'h000;
    rom[3925 ] = 12'h000;
    rom[3926 ] = 12'h000;
    rom[3927 ] = 12'h000;
    rom[3928 ] = 12'h000;
    rom[3929 ] = 12'h000;
    rom[3930 ] = 12'h000;
    rom[3931 ] = 12'h000;
    rom[3932 ] = 12'h000;
    rom[3933 ] = 12'h000;
    rom[3934 ] = 12'h000;
    rom[3935 ] = 12'h000;
    rom[3936 ] = 12'h000;
    rom[3937 ] = 12'h000;
    rom[3938 ] = 12'h000;
    rom[3939 ] = 12'h000;
    rom[3940 ] = 12'h000;
    rom[3941 ] = 12'h000;
    rom[3942 ] = 12'h000;
    rom[3943 ] = 12'h000;
    rom[3944 ] = 12'h000;
    rom[3945 ] = 12'h000;
    rom[3946 ] = 12'h000;
    rom[3947 ] = 12'h3a2;
    rom[3948 ] = 12'h3a2;
    rom[3949 ] = 12'h3a2;
    rom[3950 ] = 12'h3a2;
    rom[3951 ] = 12'h3a2;
    rom[3952 ] = 12'h3a2;
    rom[3953 ] = 12'h3a2;
    rom[3954 ] = 12'h3a2;
    rom[3955 ] = 12'h3a2;
    rom[3956 ] = 12'h3a2;
    rom[3957 ] = 12'h3a2;
    rom[3958 ] = 12'h0f0;
    rom[3959 ] = 12'h000;
    rom[3960 ] = 12'h000;
    rom[3961 ] = 12'h000;
    rom[3962 ] = 12'h000;
    rom[3963 ] = 12'h000;
    rom[3964 ] = 12'h000;
    rom[3965 ] = 12'h000;
    rom[3966 ] = 12'h000;
    rom[3967 ] = 12'h000;
    rom[3968 ] = 12'h000;
    rom[3969 ] = 12'h000;
    rom[3970 ] = 12'h000;
    rom[3971 ] = 12'h000;
    rom[3972 ] = 12'h000;
    rom[3973 ] = 12'h000;
    rom[3974 ] = 12'h000;
    rom[3975 ] = 12'h000;
    rom[3976 ] = 12'h000;
    rom[3977 ] = 12'hbb3;
    rom[3978 ] = 12'hbb3;
    rom[3979 ] = 12'hbb3;
    rom[3980 ] = 12'hbb3;
    rom[3981 ] = 12'hbb3;
    rom[3982 ] = 12'hbb3;
    rom[3983 ] = 12'hbb2;
    rom[3984 ] = 12'hbb2;
    rom[3985 ] = 12'hca2;
    rom[3986 ] = 12'hca2;
    rom[3987 ] = 12'hca2;
    rom[3988 ] = 12'hca2;
    rom[3989 ] = 12'hca2;
    rom[3990 ] = 12'hca2;
    rom[3991 ] = 12'hca2;
    rom[3992 ] = 12'hca2;
    rom[3993 ] = 12'hca2;
    rom[3994 ] = 12'hca1;
    rom[3995 ] = 12'h000;
    rom[3996 ] = 12'h000;
    rom[3997 ] = 12'h000;
    rom[3998 ] = 12'h000;
    rom[3999 ] = 12'h000;
    rom[4000 ] = 12'h000;
    rom[4001 ] = 12'h000;
    rom[4002 ] = 12'h000;
    rom[4003 ] = 12'h000;
    rom[4004 ] = 12'h000;
    rom[4005 ] = 12'h000;
    rom[4006 ] = 12'h000;
    rom[4007 ] = 12'h000;
    rom[4008 ] = 12'h000;
    rom[4009 ] = 12'h000;
    rom[4010 ] = 12'h000;
    rom[4011 ] = 12'h000;
    rom[4012 ] = 12'h000;
    rom[4013 ] = 12'h000;
    rom[4014 ] = 12'h000;
    rom[4015 ] = 12'h000;
    rom[4016 ] = 12'h000;
    rom[4017 ] = 12'h000;
    rom[4018 ] = 12'h000;
    rom[4019 ] = 12'h000;
    rom[4020 ] = 12'h000;
    rom[4021 ] = 12'h000;
    rom[4022 ] = 12'h000;
    rom[4023 ] = 12'h000;
    rom[4024 ] = 12'h000;
    rom[4025 ] = 12'h000;
    rom[4026 ] = 12'h000;
    rom[4027 ] = 12'h000;
    rom[4028 ] = 12'h000;
    rom[4029 ] = 12'h000;
    rom[4030 ] = 12'h000;
    rom[4031 ] = 12'h000;
    rom[4032 ] = 12'h000;
    rom[4033 ] = 12'h000;
    rom[4034 ] = 12'h000;
    rom[4035 ] = 12'h000;
    rom[4036 ] = 12'h000;
    rom[4037 ] = 12'h000;
    rom[4038 ] = 12'h000;
    rom[4039 ] = 12'h000;
    rom[4040 ] = 12'h000;
    rom[4041 ] = 12'h000;
    rom[4042 ] = 12'h000;
    rom[4043 ] = 12'h000;
    rom[4044 ] = 12'h000;
    rom[4045 ] = 12'h000;
    rom[4046 ] = 12'h000;
    rom[4047 ] = 12'h000;
    rom[4048 ] = 12'h000;
    rom[4049 ] = 12'h000;
    rom[4050 ] = 12'h000;
    rom[4051 ] = 12'h000;
    rom[4052 ] = 12'h000;
    rom[4053 ] = 12'h000;
    rom[4054 ] = 12'h000;
    rom[4055 ] = 12'h000;
    rom[4056 ] = 12'h000;
    rom[4057 ] = 12'h000;
    rom[4058 ] = 12'h000;
    rom[4059 ] = 12'h000;
    rom[4060 ] = 12'h000;
    rom[4061 ] = 12'h000;
    rom[4062 ] = 12'h000;
    rom[4063 ] = 12'h000;
    rom[4064 ] = 12'h000;
    rom[4065 ] = 12'h000;
    rom[4066 ] = 12'h000;
    rom[4067 ] = 12'h000;
    rom[4068 ] = 12'h000;
    rom[4069 ] = 12'h000;
    rom[4070 ] = 12'h000;
    rom[4071 ] = 12'h000;
    rom[4072 ] = 12'h000;
    rom[4073 ] = 12'h000;
    rom[4074 ] = 12'h3a2;
    rom[4075 ] = 12'h3a2;
    rom[4076 ] = 12'h3a2;
    rom[4077 ] = 12'h3a2;
    rom[4078 ] = 12'h3a2;
    rom[4079 ] = 12'h3a2;
    rom[4080 ] = 12'h3a2;
    rom[4081 ] = 12'h3a2;
    rom[4082 ] = 12'h3a2;
    rom[4083 ] = 12'h3a2;
    rom[4084 ] = 12'h3a2;
    rom[4085 ] = 12'h3a2;
    rom[4086 ] = 12'h3a2;
    rom[4087 ] = 12'h000;
    rom[4088 ] = 12'h000;
    rom[4089 ] = 12'h000;
    rom[4090 ] = 12'h000;
    rom[4091 ] = 12'h000;
    rom[4092 ] = 12'h000;
    rom[4093 ] = 12'h000;
    rom[4094 ] = 12'h000;
    rom[4095 ] = 12'h000;
    rom[4096 ] = 12'h000;
    rom[4097 ] = 12'h000;
    rom[4098 ] = 12'h000;
    rom[4099 ] = 12'h000;
    rom[4100 ] = 12'h000;
    rom[4101 ] = 12'h000;
    rom[4102 ] = 12'h000;
    rom[4103 ] = 12'h000;
    rom[4104 ] = 12'hab3;
    rom[4105 ] = 12'hbb3;
    rom[4106 ] = 12'hbb3;
    rom[4107 ] = 12'hbb3;
    rom[4108 ] = 12'hbb3;
    rom[4109 ] = 12'hbb3;
    rom[4110 ] = 12'hbb3;
    rom[4111 ] = 12'hbb3;
    rom[4112 ] = 12'hbb3;
    rom[4113 ] = 12'hbb2;
    rom[4114 ] = 12'hbb2;
    rom[4115 ] = 12'hba2;
    rom[4116 ] = 12'hca2;
    rom[4117 ] = 12'hca2;
    rom[4118 ] = 12'hca2;
    rom[4119 ] = 12'hca2;
    rom[4120 ] = 12'hca2;
    rom[4121 ] = 12'hca2;
    rom[4122 ] = 12'h000;
    rom[4123 ] = 12'h000;
    rom[4124 ] = 12'h000;
    rom[4125 ] = 12'h000;
    rom[4126 ] = 12'h000;
    rom[4127 ] = 12'h000;
    rom[4128 ] = 12'h000;
    rom[4129 ] = 12'h000;
    rom[4130 ] = 12'h000;
    rom[4131 ] = 12'h000;
    rom[4132 ] = 12'h000;
    rom[4133 ] = 12'h000;
    rom[4134 ] = 12'h000;
    rom[4135 ] = 12'h000;
    rom[4136 ] = 12'h000;
    rom[4137 ] = 12'h000;
    rom[4138 ] = 12'h000;
    rom[4139 ] = 12'h000;
    rom[4140 ] = 12'h000;
    rom[4141 ] = 12'h000;
    rom[4142 ] = 12'h000;
    rom[4143 ] = 12'h000;
    rom[4144 ] = 12'h000;
    rom[4145 ] = 12'h000;
    rom[4146 ] = 12'h000;
    rom[4147 ] = 12'h000;
    rom[4148 ] = 12'h000;
    rom[4149 ] = 12'h000;
    rom[4150 ] = 12'h000;
    rom[4151 ] = 12'h000;
    rom[4152 ] = 12'h000;
    rom[4153 ] = 12'h000;
    rom[4154 ] = 12'h000;
    rom[4155 ] = 12'h000;
    rom[4156 ] = 12'h000;
    rom[4157 ] = 12'h000;
    rom[4158 ] = 12'h000;
    rom[4159 ] = 12'h000;
    rom[4160 ] = 12'h000;
    rom[4161 ] = 12'h000;
    rom[4162 ] = 12'h000;
    rom[4163 ] = 12'h000;
    rom[4164 ] = 12'h000;
    rom[4165 ] = 12'h000;
    rom[4166 ] = 12'h000;
    rom[4167 ] = 12'h000;
    rom[4168 ] = 12'h000;
    rom[4169 ] = 12'h000;
    rom[4170 ] = 12'h000;
    rom[4171 ] = 12'h000;
    rom[4172 ] = 12'h000;
    rom[4173 ] = 12'h000;
    rom[4174 ] = 12'h000;
    rom[4175 ] = 12'h000;
    rom[4176 ] = 12'h000;
    rom[4177 ] = 12'h000;
    rom[4178 ] = 12'h000;
    rom[4179 ] = 12'h000;
    rom[4180 ] = 12'h000;
    rom[4181 ] = 12'h000;
    rom[4182 ] = 12'h000;
    rom[4183 ] = 12'h000;
    rom[4184 ] = 12'h000;
    rom[4185 ] = 12'h000;
    rom[4186 ] = 12'h000;
    rom[4187 ] = 12'h000;
    rom[4188 ] = 12'h000;
    rom[4189 ] = 12'h000;
    rom[4190 ] = 12'h000;
    rom[4191 ] = 12'h000;
    rom[4192 ] = 12'h000;
    rom[4193 ] = 12'h000;
    rom[4194 ] = 12'h000;
    rom[4195 ] = 12'h000;
    rom[4196 ] = 12'h000;
    rom[4197 ] = 12'h000;
    rom[4198 ] = 12'h000;
    rom[4199 ] = 12'h000;
    rom[4200 ] = 12'h3a2;
    rom[4201 ] = 12'h3a2;
    rom[4202 ] = 12'h3a2;
    rom[4203 ] = 12'h3a2;
    rom[4204 ] = 12'h3a2;
    rom[4205 ] = 12'h3a2;
    rom[4206 ] = 12'h3a2;
    rom[4207 ] = 12'h3a2;
    rom[4208 ] = 12'h3a2;
    rom[4209 ] = 12'h3a2;
    rom[4210 ] = 12'h3a2;
    rom[4211 ] = 12'h3a2;
    rom[4212 ] = 12'h3a2;
    rom[4213 ] = 12'h3a2;
    rom[4214 ] = 12'h3a2;
    rom[4215 ] = 12'h3a2;
    rom[4216 ] = 12'h000;
    rom[4217 ] = 12'h000;
    rom[4218 ] = 12'h000;
    rom[4219 ] = 12'h000;
    rom[4220 ] = 12'h000;
    rom[4221 ] = 12'h000;
    rom[4222 ] = 12'h000;
    rom[4223 ] = 12'h000;
    rom[4224 ] = 12'h000;
    rom[4225 ] = 12'h000;
    rom[4226 ] = 12'h000;
    rom[4227 ] = 12'h000;
    rom[4228 ] = 12'h000;
    rom[4229 ] = 12'h000;
    rom[4230 ] = 12'h000;
    rom[4231 ] = 12'h000;
    rom[4232 ] = 12'hab3;
    rom[4233 ] = 12'hab3;
    rom[4234 ] = 12'hab3;
    rom[4235 ] = 12'hab3;
    rom[4236 ] = 12'hbb3;
    rom[4237 ] = 12'hbb3;
    rom[4238 ] = 12'hbb3;
    rom[4239 ] = 12'hbb3;
    rom[4240 ] = 12'hbb3;
    rom[4241 ] = 12'hbb3;
    rom[4242 ] = 12'hbb3;
    rom[4243 ] = 12'hbb3;
    rom[4244 ] = 12'hbb2;
    rom[4245 ] = 12'hbb2;
    rom[4246 ] = 12'hca2;
    rom[4247 ] = 12'hca2;
    rom[4248 ] = 12'hca2;
    rom[4249 ] = 12'hca2;
    rom[4250 ] = 12'h000;
    rom[4251 ] = 12'h000;
    rom[4252 ] = 12'h000;
    rom[4253 ] = 12'h000;
    rom[4254 ] = 12'h000;
    rom[4255 ] = 12'h000;
    rom[4256 ] = 12'h000;
    rom[4257 ] = 12'h000;
    rom[4258 ] = 12'h000;
    rom[4259 ] = 12'h000;
    rom[4260 ] = 12'h000;
    rom[4261 ] = 12'h000;
    rom[4262 ] = 12'h000;
    rom[4263 ] = 12'h000;
    rom[4264 ] = 12'h000;
    rom[4265 ] = 12'h000;
    rom[4266 ] = 12'h000;
    rom[4267 ] = 12'h000;
    rom[4268 ] = 12'h000;
    rom[4269 ] = 12'h000;
    rom[4270 ] = 12'h000;
    rom[4271 ] = 12'h000;
    rom[4272 ] = 12'h000;
    rom[4273 ] = 12'h000;
    rom[4274 ] = 12'h000;
    rom[4275 ] = 12'h000;
    rom[4276 ] = 12'h000;
    rom[4277 ] = 12'h000;
    rom[4278 ] = 12'h000;
    rom[4279 ] = 12'h000;
    rom[4280 ] = 12'h000;
    rom[4281 ] = 12'h000;
    rom[4282 ] = 12'h000;
    rom[4283 ] = 12'h000;
    rom[4284 ] = 12'h000;
    rom[4285 ] = 12'h000;
    rom[4286 ] = 12'h000;
    rom[4287 ] = 12'h000;
    rom[4288 ] = 12'h000;
    rom[4289 ] = 12'h000;
    rom[4290 ] = 12'h000;
    rom[4291 ] = 12'h000;
    rom[4292 ] = 12'h000;
    rom[4293 ] = 12'h000;
    rom[4294 ] = 12'h000;
    rom[4295 ] = 12'h000;
    rom[4296 ] = 12'h000;
    rom[4297 ] = 12'h000;
    rom[4298 ] = 12'h000;
    rom[4299 ] = 12'h000;
    rom[4300 ] = 12'h000;
    rom[4301 ] = 12'h000;
    rom[4302 ] = 12'h000;
    rom[4303 ] = 12'h000;
    rom[4304 ] = 12'h000;
    rom[4305 ] = 12'h000;
    rom[4306 ] = 12'h000;
    rom[4307 ] = 12'h000;
    rom[4308 ] = 12'h000;
    rom[4309 ] = 12'h000;
    rom[4310 ] = 12'h000;
    rom[4311 ] = 12'h000;
    rom[4312 ] = 12'h000;
    rom[4313 ] = 12'h000;
    rom[4314 ] = 12'h000;
    rom[4315 ] = 12'h000;
    rom[4316 ] = 12'h000;
    rom[4317 ] = 12'h000;
    rom[4318 ] = 12'h000;
    rom[4319 ] = 12'h000;
    rom[4320 ] = 12'h000;
    rom[4321 ] = 12'h000;
    rom[4322 ] = 12'h000;
    rom[4323 ] = 12'h000;
    rom[4324 ] = 12'h000;
    rom[4325 ] = 12'h000;
    rom[4326 ] = 12'h000;
    rom[4327 ] = 12'h3a2;
    rom[4328 ] = 12'h3a2;
    rom[4329 ] = 12'h3a2;
    rom[4330 ] = 12'h3a2;
    rom[4331 ] = 12'h3a2;
    rom[4332 ] = 12'h3a2;
    rom[4333 ] = 12'h3a2;
    rom[4334 ] = 12'h3a2;
    rom[4335 ] = 12'h3a2;
    rom[4336 ] = 12'h3a2;
    rom[4337 ] = 12'h3a2;
    rom[4338 ] = 12'h3a2;
    rom[4339 ] = 12'h3a2;
    rom[4340 ] = 12'h3a2;
    rom[4341 ] = 12'h3a2;
    rom[4342 ] = 12'h3a2;
    rom[4343 ] = 12'h3a2;
    rom[4344 ] = 12'h000;
    rom[4345 ] = 12'h000;
    rom[4346 ] = 12'h000;
    rom[4347 ] = 12'h000;
    rom[4348 ] = 12'h000;
    rom[4349 ] = 12'h000;
    rom[4350 ] = 12'h000;
    rom[4351 ] = 12'h000;
    rom[4352 ] = 12'h000;
    rom[4353 ] = 12'h000;
    rom[4354 ] = 12'h000;
    rom[4355 ] = 12'h000;
    rom[4356 ] = 12'h000;
    rom[4357 ] = 12'h000;
    rom[4358 ] = 12'h000;
    rom[4359 ] = 12'hab4;
    rom[4360 ] = 12'hab4;
    rom[4361 ] = 12'hab4;
    rom[4362 ] = 12'hab4;
    rom[4363 ] = 12'hab3;
    rom[4364 ] = 12'hab3;
    rom[4365 ] = 12'hab3;
    rom[4366 ] = 12'hab3;
    rom[4367 ] = 12'hbb3;
    rom[4368 ] = 12'hbb3;
    rom[4369 ] = 12'hbb3;
    rom[4370 ] = 12'hbb3;
    rom[4371 ] = 12'hbb3;
    rom[4372 ] = 12'hbb3;
    rom[4373 ] = 12'hbb3;
    rom[4374 ] = 12'hbb2;
    rom[4375 ] = 12'hbb2;
    rom[4376 ] = 12'hba2;
    rom[4377 ] = 12'h000;
    rom[4378 ] = 12'h000;
    rom[4379 ] = 12'h000;
    rom[4380 ] = 12'h000;
    rom[4381 ] = 12'h000;
    rom[4382 ] = 12'h000;
    rom[4383 ] = 12'h000;
    rom[4384 ] = 12'h000;
    rom[4385 ] = 12'h000;
    rom[4386 ] = 12'h000;
    rom[4387 ] = 12'h000;
    rom[4388 ] = 12'h000;
    rom[4389 ] = 12'h000;
    rom[4390 ] = 12'h000;
    rom[4391 ] = 12'h000;
    rom[4392 ] = 12'h000;
    rom[4393 ] = 12'h000;
    rom[4394 ] = 12'h000;
    rom[4395 ] = 12'h000;
    rom[4396 ] = 12'h000;
    rom[4397 ] = 12'h000;
    rom[4398 ] = 12'h000;
    rom[4399 ] = 12'h000;
    rom[4400 ] = 12'h000;
    rom[4401 ] = 12'h000;
    rom[4402 ] = 12'h000;
    rom[4403 ] = 12'h000;
    rom[4404 ] = 12'h000;
    rom[4405 ] = 12'h000;
    rom[4406 ] = 12'h000;
    rom[4407 ] = 12'h000;
    rom[4408 ] = 12'h000;
    rom[4409 ] = 12'h000;
    rom[4410 ] = 12'h000;
    rom[4411 ] = 12'h000;
    rom[4412 ] = 12'h000;
    rom[4413 ] = 12'h000;
    rom[4414 ] = 12'h000;
    rom[4415 ] = 12'h000;
    rom[4416 ] = 12'h000;
    rom[4417 ] = 12'h000;
    rom[4418 ] = 12'h000;
    rom[4419 ] = 12'h000;
    rom[4420 ] = 12'h000;
    rom[4421 ] = 12'h000;
    rom[4422 ] = 12'h000;
    rom[4423 ] = 12'h000;
    rom[4424 ] = 12'h000;
    rom[4425 ] = 12'h000;
    rom[4426 ] = 12'h000;
    rom[4427 ] = 12'h000;
    rom[4428 ] = 12'h000;
    rom[4429 ] = 12'h000;
    rom[4430 ] = 12'h000;
    rom[4431 ] = 12'h000;
    rom[4432 ] = 12'h000;
    rom[4433 ] = 12'h000;
    rom[4434 ] = 12'h000;
    rom[4435 ] = 12'h000;
    rom[4436 ] = 12'h000;
    rom[4437 ] = 12'h000;
    rom[4438 ] = 12'h000;
    rom[4439 ] = 12'h000;
    rom[4440 ] = 12'h000;
    rom[4441 ] = 12'h000;
    rom[4442 ] = 12'h000;
    rom[4443 ] = 12'h000;
    rom[4444 ] = 12'h000;
    rom[4445 ] = 12'h000;
    rom[4446 ] = 12'h000;
    rom[4447 ] = 12'h000;
    rom[4448 ] = 12'h000;
    rom[4449 ] = 12'h000;
    rom[4450 ] = 12'h000;
    rom[4451 ] = 12'h000;
    rom[4452 ] = 12'h000;
    rom[4453 ] = 12'h4a1;
    rom[4454 ] = 12'h3a2;
    rom[4455 ] = 12'h3a2;
    rom[4456 ] = 12'h3a2;
    rom[4457 ] = 12'h3a2;
    rom[4458 ] = 12'h3a2;
    rom[4459 ] = 12'h3a2;
    rom[4460 ] = 12'h3a2;
    rom[4461 ] = 12'h3a2;
    rom[4462 ] = 12'h3a2;
    rom[4463 ] = 12'h3a2;
    rom[4464 ] = 12'h3a2;
    rom[4465 ] = 12'h3a2;
    rom[4466 ] = 12'h3a2;
    rom[4467 ] = 12'h3a2;
    rom[4468 ] = 12'h3a2;
    rom[4469 ] = 12'h3a2;
    rom[4470 ] = 12'h3a2;
    rom[4471 ] = 12'h3a2;
    rom[4472 ] = 12'h3a2;
    rom[4473 ] = 12'h000;
    rom[4474 ] = 12'h000;
    rom[4475 ] = 12'h000;
    rom[4476 ] = 12'h000;
    rom[4477 ] = 12'h000;
    rom[4478 ] = 12'h000;
    rom[4479 ] = 12'h000;
    rom[4480 ] = 12'h000;
    rom[4481 ] = 12'h000;
    rom[4482 ] = 12'h000;
    rom[4483 ] = 12'h000;
    rom[4484 ] = 12'h000;
    rom[4485 ] = 12'h000;
    rom[4486 ] = 12'h000;
    rom[4487 ] = 12'hab4;
    rom[4488 ] = 12'hab4;
    rom[4489 ] = 12'hab4;
    rom[4490 ] = 12'hab4;
    rom[4491 ] = 12'hab4;
    rom[4492 ] = 12'hab4;
    rom[4493 ] = 12'hab3;
    rom[4494 ] = 12'hab3;
    rom[4495 ] = 12'hab3;
    rom[4496 ] = 12'hab3;
    rom[4497 ] = 12'hbb3;
    rom[4498 ] = 12'hbb3;
    rom[4499 ] = 12'hbb3;
    rom[4500 ] = 12'hbb3;
    rom[4501 ] = 12'hbb3;
    rom[4502 ] = 12'hbb3;
    rom[4503 ] = 12'hbb3;
    rom[4504 ] = 12'h000;
    rom[4505 ] = 12'h000;
    rom[4506 ] = 12'h000;
    rom[4507 ] = 12'h000;
    rom[4508 ] = 12'h000;
    rom[4509 ] = 12'h000;
    rom[4510 ] = 12'h000;
    rom[4511 ] = 12'h000;
    rom[4512 ] = 12'h000;
    rom[4513 ] = 12'h000;
    rom[4514 ] = 12'h000;
    rom[4515 ] = 12'h000;
    rom[4516 ] = 12'h000;
    rom[4517 ] = 12'h000;
    rom[4518 ] = 12'h000;
    rom[4519 ] = 12'h000;
    rom[4520 ] = 12'h000;
    rom[4521 ] = 12'h000;
    rom[4522 ] = 12'h000;
    rom[4523 ] = 12'h000;
    rom[4524 ] = 12'h000;
    rom[4525 ] = 12'h000;
    rom[4526 ] = 12'h000;
    rom[4527 ] = 12'h000;
    rom[4528 ] = 12'h000;
    rom[4529 ] = 12'h000;
    rom[4530 ] = 12'h000;
    rom[4531 ] = 12'h000;
    rom[4532 ] = 12'h000;
    rom[4533 ] = 12'h000;
    rom[4534 ] = 12'h000;
    rom[4535 ] = 12'h000;
    rom[4536 ] = 12'h000;
    rom[4537 ] = 12'h000;
    rom[4538 ] = 12'h000;
    rom[4539 ] = 12'h000;
    rom[4540 ] = 12'h000;
    rom[4541 ] = 12'h000;
    rom[4542 ] = 12'h000;
    rom[4543 ] = 12'h000;
    rom[4544 ] = 12'h000;
    rom[4545 ] = 12'h000;
    rom[4546 ] = 12'h000;
    rom[4547 ] = 12'h000;
    rom[4548 ] = 12'h000;
    rom[4549 ] = 12'h000;
    rom[4550 ] = 12'h000;
    rom[4551 ] = 12'h000;
    rom[4552 ] = 12'h000;
    rom[4553 ] = 12'h000;
    rom[4554 ] = 12'h000;
    rom[4555 ] = 12'h000;
    rom[4556 ] = 12'h000;
    rom[4557 ] = 12'h000;
    rom[4558 ] = 12'h000;
    rom[4559 ] = 12'h000;
    rom[4560 ] = 12'h000;
    rom[4561 ] = 12'h000;
    rom[4562 ] = 12'h000;
    rom[4563 ] = 12'h000;
    rom[4564 ] = 12'h000;
    rom[4565 ] = 12'h000;
    rom[4566 ] = 12'h000;
    rom[4567 ] = 12'h000;
    rom[4568 ] = 12'h000;
    rom[4569 ] = 12'h000;
    rom[4570 ] = 12'h000;
    rom[4571 ] = 12'h000;
    rom[4572 ] = 12'h000;
    rom[4573 ] = 12'h000;
    rom[4574 ] = 12'h000;
    rom[4575 ] = 12'h000;
    rom[4576 ] = 12'h000;
    rom[4577 ] = 12'h000;
    rom[4578 ] = 12'h000;
    rom[4579 ] = 12'h000;
    rom[4580 ] = 12'h3a2;
    rom[4581 ] = 12'h3a2;
    rom[4582 ] = 12'h3a2;
    rom[4583 ] = 12'h3a2;
    rom[4584 ] = 12'h3a2;
    rom[4585 ] = 12'h3a2;
    rom[4586 ] = 12'h3a2;
    rom[4587 ] = 12'h3a2;
    rom[4588 ] = 12'h3a2;
    rom[4589 ] = 12'h3a2;
    rom[4590 ] = 12'h3a2;
    rom[4591 ] = 12'h3a2;
    rom[4592 ] = 12'h3a2;
    rom[4593 ] = 12'h3a2;
    rom[4594 ] = 12'h3a2;
    rom[4595 ] = 12'h3a2;
    rom[4596 ] = 12'h3a2;
    rom[4597 ] = 12'h3a2;
    rom[4598 ] = 12'h3a2;
    rom[4599 ] = 12'h3a2;
    rom[4600 ] = 12'h3a2;
    rom[4601 ] = 12'h000;
    rom[4602 ] = 12'h000;
    rom[4603 ] = 12'h000;
    rom[4604 ] = 12'h000;
    rom[4605 ] = 12'h000;
    rom[4606 ] = 12'h000;
    rom[4607 ] = 12'h000;
    rom[4608 ] = 12'h000;
    rom[4609 ] = 12'h000;
    rom[4610 ] = 12'h000;
    rom[4611 ] = 12'h000;
    rom[4612 ] = 12'h000;
    rom[4613 ] = 12'h000;
    rom[4614 ] = 12'h9b4;
    rom[4615 ] = 12'h9b4;
    rom[4616 ] = 12'h9b4;
    rom[4617 ] = 12'h9b4;
    rom[4618 ] = 12'hab4;
    rom[4619 ] = 12'hab4;
    rom[4620 ] = 12'hab4;
    rom[4621 ] = 12'hab4;
    rom[4622 ] = 12'hab4;
    rom[4623 ] = 12'hab4;
    rom[4624 ] = 12'hab3;
    rom[4625 ] = 12'hab3;
    rom[4626 ] = 12'hab3;
    rom[4627 ] = 12'hab3;
    rom[4628 ] = 12'hbb3;
    rom[4629 ] = 12'hbb3;
    rom[4630 ] = 12'hbb3;
    rom[4631 ] = 12'h000;
    rom[4632 ] = 12'h000;
    rom[4633 ] = 12'h000;
    rom[4634 ] = 12'h000;
    rom[4635 ] = 12'h000;
    rom[4636 ] = 12'h000;
    rom[4637 ] = 12'h000;
    rom[4638 ] = 12'h000;
    rom[4639 ] = 12'h000;
    rom[4640 ] = 12'h000;
    rom[4641 ] = 12'h000;
    rom[4642 ] = 12'h000;
    rom[4643 ] = 12'h000;
    rom[4644 ] = 12'h000;
    rom[4645 ] = 12'h000;
    rom[4646 ] = 12'h000;
    rom[4647 ] = 12'h000;
    rom[4648 ] = 12'h000;
    rom[4649 ] = 12'h000;
    rom[4650 ] = 12'h000;
    rom[4651 ] = 12'h000;
    rom[4652 ] = 12'h000;
    rom[4653 ] = 12'h000;
    rom[4654 ] = 12'h000;
    rom[4655 ] = 12'h000;
    rom[4656 ] = 12'h000;
    rom[4657 ] = 12'h000;
    rom[4658 ] = 12'h000;
    rom[4659 ] = 12'h000;
    rom[4660 ] = 12'h000;
    rom[4661 ] = 12'h000;
    rom[4662 ] = 12'h000;
    rom[4663 ] = 12'h000;
    rom[4664 ] = 12'h000;
    rom[4665 ] = 12'h000;
    rom[4666 ] = 12'h000;
    rom[4667 ] = 12'h000;
    rom[4668 ] = 12'h000;
    rom[4669 ] = 12'h000;
    rom[4670 ] = 12'h000;
    rom[4671 ] = 12'h000;
    rom[4672 ] = 12'h000;
    rom[4673 ] = 12'h000;
    rom[4674 ] = 12'h000;
    rom[4675 ] = 12'h000;
    rom[4676 ] = 12'h000;
    rom[4677 ] = 12'h000;
    rom[4678 ] = 12'h000;
    rom[4679 ] = 12'h000;
    rom[4680 ] = 12'h000;
    rom[4681 ] = 12'h000;
    rom[4682 ] = 12'h000;
    rom[4683 ] = 12'h000;
    rom[4684 ] = 12'h000;
    rom[4685 ] = 12'h000;
    rom[4686 ] = 12'h000;
    rom[4687 ] = 12'h000;
    rom[4688 ] = 12'h000;
    rom[4689 ] = 12'h000;
    rom[4690 ] = 12'h000;
    rom[4691 ] = 12'h000;
    rom[4692 ] = 12'h000;
    rom[4693 ] = 12'h000;
    rom[4694 ] = 12'h000;
    rom[4695 ] = 12'h000;
    rom[4696 ] = 12'h000;
    rom[4697 ] = 12'h000;
    rom[4698 ] = 12'h000;
    rom[4699 ] = 12'h000;
    rom[4700 ] = 12'h000;
    rom[4701 ] = 12'h000;
    rom[4702 ] = 12'h000;
    rom[4703 ] = 12'h000;
    rom[4704 ] = 12'h000;
    rom[4705 ] = 12'h000;
    rom[4706 ] = 12'h000;
    rom[4707 ] = 12'h3a2;
    rom[4708 ] = 12'h3a2;
    rom[4709 ] = 12'h3a2;
    rom[4710 ] = 12'h3a2;
    rom[4711 ] = 12'h3a2;
    rom[4712 ] = 12'h3a2;
    rom[4713 ] = 12'h3a2;
    rom[4714 ] = 12'h3a2;
    rom[4715 ] = 12'h3a2;
    rom[4716 ] = 12'h3a2;
    rom[4717 ] = 12'h3a2;
    rom[4718 ] = 12'h3a2;
    rom[4719 ] = 12'h3a2;
    rom[4720 ] = 12'h3a2;
    rom[4721 ] = 12'h3a2;
    rom[4722 ] = 12'h3a2;
    rom[4723 ] = 12'h3a2;
    rom[4724 ] = 12'h3a2;
    rom[4725 ] = 12'h3a2;
    rom[4726 ] = 12'h3a2;
    rom[4727 ] = 12'h3a2;
    rom[4728 ] = 12'h3a2;
    rom[4729 ] = 12'h3a2;
    rom[4730 ] = 12'h000;
    rom[4731 ] = 12'h000;
    rom[4732 ] = 12'h000;
    rom[4733 ] = 12'h000;
    rom[4734 ] = 12'h000;
    rom[4735 ] = 12'h000;
    rom[4736 ] = 12'h000;
    rom[4737 ] = 12'h000;
    rom[4738 ] = 12'h000;
    rom[4739 ] = 12'h000;
    rom[4740 ] = 12'h000;
    rom[4741 ] = 12'h000;
    rom[4742 ] = 12'h9b4;
    rom[4743 ] = 12'h9b4;
    rom[4744 ] = 12'h9b4;
    rom[4745 ] = 12'h9b4;
    rom[4746 ] = 12'h9b4;
    rom[4747 ] = 12'h9b4;
    rom[4748 ] = 12'hab4;
    rom[4749 ] = 12'hab4;
    rom[4750 ] = 12'hab4;
    rom[4751 ] = 12'hab4;
    rom[4752 ] = 12'hab4;
    rom[4753 ] = 12'hab4;
    rom[4754 ] = 12'hab3;
    rom[4755 ] = 12'hab3;
    rom[4756 ] = 12'hab3;
    rom[4757 ] = 12'hab3;
    rom[4758 ] = 12'hbb3;
    rom[4759 ] = 12'h000;
    rom[4760 ] = 12'h000;
    rom[4761 ] = 12'h000;
    rom[4762 ] = 12'h000;
    rom[4763 ] = 12'h000;
    rom[4764 ] = 12'h000;
    rom[4765 ] = 12'h000;
    rom[4766 ] = 12'h000;
    rom[4767 ] = 12'h000;
    rom[4768 ] = 12'h000;
    rom[4769 ] = 12'h000;
    rom[4770 ] = 12'h000;
    rom[4771 ] = 12'h000;
    rom[4772 ] = 12'h000;
    rom[4773 ] = 12'h000;
    rom[4774 ] = 12'h000;
    rom[4775 ] = 12'h000;
    rom[4776 ] = 12'h000;
    rom[4777 ] = 12'h000;
    rom[4778 ] = 12'h000;
    rom[4779 ] = 12'h000;
    rom[4780 ] = 12'h000;
    rom[4781 ] = 12'h000;
    rom[4782 ] = 12'h000;
    rom[4783 ] = 12'h000;
    rom[4784 ] = 12'h000;
    rom[4785 ] = 12'h000;
    rom[4786 ] = 12'h000;
    rom[4787 ] = 12'h000;
    rom[4788 ] = 12'h000;
    rom[4789 ] = 12'h000;
    rom[4790 ] = 12'h000;
    rom[4791 ] = 12'h000;
    rom[4792 ] = 12'h000;
    rom[4793 ] = 12'h000;
    rom[4794 ] = 12'h000;
    rom[4795 ] = 12'h000;
    rom[4796 ] = 12'h000;
    rom[4797 ] = 12'h000;
    rom[4798 ] = 12'h000;
    rom[4799 ] = 12'h000;
    rom[4800 ] = 12'h000;
    rom[4801 ] = 12'h000;
    rom[4802 ] = 12'h000;
    rom[4803 ] = 12'h000;
    rom[4804 ] = 12'h000;
    rom[4805 ] = 12'h000;
    rom[4806 ] = 12'h000;
    rom[4807 ] = 12'h000;
    rom[4808 ] = 12'h000;
    rom[4809 ] = 12'h000;
    rom[4810 ] = 12'h000;
    rom[4811 ] = 12'h000;
    rom[4812 ] = 12'h000;
    rom[4813 ] = 12'h000;
    rom[4814 ] = 12'h000;
    rom[4815 ] = 12'h000;
    rom[4816 ] = 12'h000;
    rom[4817 ] = 12'h000;
    rom[4818 ] = 12'h000;
    rom[4819 ] = 12'h000;
    rom[4820 ] = 12'h000;
    rom[4821 ] = 12'h000;
    rom[4822 ] = 12'h000;
    rom[4823 ] = 12'h000;
    rom[4824 ] = 12'h000;
    rom[4825 ] = 12'h000;
    rom[4826 ] = 12'h000;
    rom[4827 ] = 12'h000;
    rom[4828 ] = 12'h000;
    rom[4829 ] = 12'h000;
    rom[4830 ] = 12'h000;
    rom[4831 ] = 12'h000;
    rom[4832 ] = 12'h000;
    rom[4833 ] = 12'h392;
    rom[4834 ] = 12'h3a2;
    rom[4835 ] = 12'h3a2;
    rom[4836 ] = 12'h3a2;
    rom[4837 ] = 12'h3a2;
    rom[4838 ] = 12'h3a2;
    rom[4839 ] = 12'h3a2;
    rom[4840 ] = 12'h3a2;
    rom[4841 ] = 12'h3a2;
    rom[4842 ] = 12'h3a2;
    rom[4843 ] = 12'h3a2;
    rom[4844 ] = 12'h3a2;
    rom[4845 ] = 12'h3a2;
    rom[4846 ] = 12'h3a2;
    rom[4847 ] = 12'h3a2;
    rom[4848 ] = 12'h3a2;
    rom[4849 ] = 12'h3a2;
    rom[4850 ] = 12'h3a2;
    rom[4851 ] = 12'h3a2;
    rom[4852 ] = 12'h3a2;
    rom[4853 ] = 12'h3a2;
    rom[4854 ] = 12'h3a2;
    rom[4855 ] = 12'h3a2;
    rom[4856 ] = 12'h3a2;
    rom[4857 ] = 12'h3a2;
    rom[4858 ] = 12'h000;
    rom[4859 ] = 12'h000;
    rom[4860 ] = 12'h000;
    rom[4861 ] = 12'h000;
    rom[4862 ] = 12'h000;
    rom[4863 ] = 12'h000;
    rom[4864 ] = 12'h000;
    rom[4865 ] = 12'h000;
    rom[4866 ] = 12'h000;
    rom[4867 ] = 12'h000;
    rom[4868 ] = 12'h000;
    rom[4869 ] = 12'h9b5;
    rom[4870 ] = 12'h9b5;
    rom[4871 ] = 12'h9b5;
    rom[4872 ] = 12'h9b5;
    rom[4873 ] = 12'h9b4;
    rom[4874 ] = 12'h9b4;
    rom[4875 ] = 12'h9b4;
    rom[4876 ] = 12'h9b4;
    rom[4877 ] = 12'h9b4;
    rom[4878 ] = 12'h9b4;
    rom[4879 ] = 12'hab4;
    rom[4880 ] = 12'hab4;
    rom[4881 ] = 12'hab4;
    rom[4882 ] = 12'hab4;
    rom[4883 ] = 12'hab4;
    rom[4884 ] = 12'hab4;
    rom[4885 ] = 12'hab3;
    rom[4886 ] = 12'h000;
    rom[4887 ] = 12'h000;
    rom[4888 ] = 12'h000;
    rom[4889 ] = 12'h000;
    rom[4890 ] = 12'h000;
    rom[4891 ] = 12'h000;
    rom[4892 ] = 12'h000;
    rom[4893 ] = 12'h000;
    rom[4894 ] = 12'h000;
    rom[4895 ] = 12'h000;
    rom[4896 ] = 12'h000;
    rom[4897 ] = 12'h000;
    rom[4898 ] = 12'h000;
    rom[4899 ] = 12'h000;
    rom[4900 ] = 12'h000;
    rom[4901 ] = 12'h000;
    rom[4902 ] = 12'h000;
    rom[4903 ] = 12'h000;
    rom[4904 ] = 12'h000;
    rom[4905 ] = 12'h000;
    rom[4906 ] = 12'h000;
    rom[4907 ] = 12'h000;
    rom[4908 ] = 12'h000;
    rom[4909 ] = 12'h000;
    rom[4910 ] = 12'h000;
    rom[4911 ] = 12'h000;
    rom[4912 ] = 12'h000;
    rom[4913 ] = 12'h000;
    rom[4914 ] = 12'h000;
    rom[4915 ] = 12'h000;
    rom[4916 ] = 12'h000;
    rom[4917 ] = 12'h000;
    rom[4918 ] = 12'h000;
    rom[4919 ] = 12'h000;
    rom[4920 ] = 12'h000;
    rom[4921 ] = 12'h000;
    rom[4922 ] = 12'h000;
    rom[4923 ] = 12'h000;
    rom[4924 ] = 12'h000;
    rom[4925 ] = 12'h000;
    rom[4926 ] = 12'h000;
    rom[4927 ] = 12'h000;
    rom[4928 ] = 12'h000;
    rom[4929 ] = 12'h000;
    rom[4930 ] = 12'h000;
    rom[4931 ] = 12'h000;
    rom[4932 ] = 12'h000;
    rom[4933 ] = 12'h000;
    rom[4934 ] = 12'h000;
    rom[4935 ] = 12'h000;
    rom[4936 ] = 12'h000;
    rom[4937 ] = 12'h000;
    rom[4938 ] = 12'h000;
    rom[4939 ] = 12'h000;
    rom[4940 ] = 12'h000;
    rom[4941 ] = 12'h000;
    rom[4942 ] = 12'h000;
    rom[4943 ] = 12'h000;
    rom[4944 ] = 12'h000;
    rom[4945 ] = 12'h000;
    rom[4946 ] = 12'h000;
    rom[4947 ] = 12'h000;
    rom[4948 ] = 12'h000;
    rom[4949 ] = 12'h000;
    rom[4950 ] = 12'h000;
    rom[4951 ] = 12'h000;
    rom[4952 ] = 12'h000;
    rom[4953 ] = 12'h000;
    rom[4954 ] = 12'h000;
    rom[4955 ] = 12'h000;
    rom[4956 ] = 12'h000;
    rom[4957 ] = 12'h000;
    rom[4958 ] = 12'h000;
    rom[4959 ] = 12'h000;
    rom[4960 ] = 12'h3a2;
    rom[4961 ] = 12'h3a2;
    rom[4962 ] = 12'h3a2;
    rom[4963 ] = 12'h3a2;
    rom[4964 ] = 12'h3a2;
    rom[4965 ] = 12'h3a2;
    rom[4966 ] = 12'h3a2;
    rom[4967 ] = 12'h3a2;
    rom[4968 ] = 12'h3a2;
    rom[4969 ] = 12'h3a2;
    rom[4970 ] = 12'h3a2;
    rom[4971 ] = 12'h3a2;
    rom[4972 ] = 12'h3a2;
    rom[4973 ] = 12'h3a2;
    rom[4974 ] = 12'h3a2;
    rom[4975 ] = 12'h3a2;
    rom[4976 ] = 12'h3a2;
    rom[4977 ] = 12'h3a2;
    rom[4978 ] = 12'h3a2;
    rom[4979 ] = 12'h3a2;
    rom[4980 ] = 12'h3a2;
    rom[4981 ] = 12'h3a2;
    rom[4982 ] = 12'h3a2;
    rom[4983 ] = 12'h3a2;
    rom[4984 ] = 12'h3a2;
    rom[4985 ] = 12'h000;
    rom[4986 ] = 12'h000;
    rom[4987 ] = 12'h000;
    rom[4988 ] = 12'h000;
    rom[4989 ] = 12'h000;
    rom[4990 ] = 12'h000;
    rom[4991 ] = 12'h000;
    rom[4992 ] = 12'h000;
    rom[4993 ] = 12'h000;
    rom[4994 ] = 12'h000;
    rom[4995 ] = 12'h000;
    rom[4996 ] = 12'h000;
    rom[4997 ] = 12'h8b5;
    rom[4998 ] = 12'h8b5;
    rom[4999 ] = 12'h9b5;
    rom[5000 ] = 12'h9b5;
    rom[5001 ] = 12'h9b5;
    rom[5002 ] = 12'h9b5;
    rom[5003 ] = 12'h9b5;
    rom[5004 ] = 12'h9b4;
    rom[5005 ] = 12'h9b4;
    rom[5006 ] = 12'h9b4;
    rom[5007 ] = 12'h9b4;
    rom[5008 ] = 12'h9b4;
    rom[5009 ] = 12'hab4;
    rom[5010 ] = 12'hab4;
    rom[5011 ] = 12'hab4;
    rom[5012 ] = 12'hab4;
    rom[5013 ] = 12'hab3;
    rom[5014 ] = 12'h000;
    rom[5015 ] = 12'h000;
    rom[5016 ] = 12'h000;
    rom[5017 ] = 12'h000;
    rom[5018 ] = 12'h000;
    rom[5019 ] = 12'h000;
    rom[5020 ] = 12'h000;
    rom[5021 ] = 12'h000;
    rom[5022 ] = 12'h000;
    rom[5023 ] = 12'h000;
    rom[5024 ] = 12'h000;
    rom[5025 ] = 12'h000;
    rom[5026 ] = 12'h000;
    rom[5027 ] = 12'h000;
    rom[5028 ] = 12'h000;
    rom[5029 ] = 12'h000;
    rom[5030 ] = 12'h000;
    rom[5031 ] = 12'h000;
    rom[5032 ] = 12'h000;
    rom[5033 ] = 12'h000;
    rom[5034 ] = 12'h000;
    rom[5035 ] = 12'h000;
    rom[5036 ] = 12'h000;
    rom[5037 ] = 12'h000;
    rom[5038 ] = 12'h000;
    rom[5039 ] = 12'h000;
    rom[5040 ] = 12'h000;
    rom[5041 ] = 12'h000;
    rom[5042 ] = 12'h000;
    rom[5043 ] = 12'h000;
    rom[5044 ] = 12'h000;
    rom[5045 ] = 12'h000;
    rom[5046 ] = 12'h000;
    rom[5047 ] = 12'h000;
    rom[5048 ] = 12'h000;
    rom[5049 ] = 12'h000;
    rom[5050 ] = 12'h000;
    rom[5051 ] = 12'h000;
    rom[5052 ] = 12'h000;
    rom[5053 ] = 12'h000;
    rom[5054 ] = 12'h000;
    rom[5055 ] = 12'h000;
    rom[5056 ] = 12'h000;
    rom[5057 ] = 12'h000;
    rom[5058 ] = 12'h000;
    rom[5059 ] = 12'h000;
    rom[5060 ] = 12'h000;
    rom[5061 ] = 12'h000;
    rom[5062 ] = 12'h000;
    rom[5063 ] = 12'h000;
    rom[5064 ] = 12'h000;
    rom[5065 ] = 12'h000;
    rom[5066 ] = 12'h000;
    rom[5067 ] = 12'h000;
    rom[5068 ] = 12'h000;
    rom[5069 ] = 12'h000;
    rom[5070 ] = 12'h000;
    rom[5071 ] = 12'h000;
    rom[5072 ] = 12'h000;
    rom[5073 ] = 12'h000;
    rom[5074 ] = 12'h000;
    rom[5075 ] = 12'h000;
    rom[5076 ] = 12'h000;
    rom[5077 ] = 12'h000;
    rom[5078 ] = 12'h000;
    rom[5079 ] = 12'h000;
    rom[5080 ] = 12'h000;
    rom[5081 ] = 12'h000;
    rom[5082 ] = 12'h000;
    rom[5083 ] = 12'h000;
    rom[5084 ] = 12'h000;
    rom[5085 ] = 12'h000;
    rom[5086 ] = 12'h000;
    rom[5087 ] = 12'h3a2;
    rom[5088 ] = 12'h3a2;
    rom[5089 ] = 12'h3a2;
    rom[5090 ] = 12'h3a2;
    rom[5091 ] = 12'h3a2;
    rom[5092 ] = 12'h3a2;
    rom[5093 ] = 12'h3a2;
    rom[5094 ] = 12'h3a2;
    rom[5095 ] = 12'h3a2;
    rom[5096 ] = 12'h3a2;
    rom[5097 ] = 12'h3a2;
    rom[5098 ] = 12'h3a2;
    rom[5099 ] = 12'h3a2;
    rom[5100 ] = 12'h3a2;
    rom[5101 ] = 12'h3a2;
    rom[5102 ] = 12'h3a2;
    rom[5103 ] = 12'h3a2;
    rom[5104 ] = 12'h3a2;
    rom[5105 ] = 12'h3a2;
    rom[5106 ] = 12'h3a2;
    rom[5107 ] = 12'h3a2;
    rom[5108 ] = 12'h3a2;
    rom[5109 ] = 12'h3a2;
    rom[5110 ] = 12'h3a2;
    rom[5111 ] = 12'h3a2;
    rom[5112 ] = 12'h000;
    rom[5113 ] = 12'h000;
    rom[5114 ] = 12'h000;
    rom[5115 ] = 12'h000;
    rom[5116 ] = 12'h000;
    rom[5117 ] = 12'h000;
    rom[5118 ] = 12'h000;
    rom[5119 ] = 12'h000;
    rom[5120 ] = 12'h000;
    rom[5121 ] = 12'h000;
    rom[5122 ] = 12'h000;
    rom[5123 ] = 12'h000;
    rom[5124 ] = 12'h8b5;
    rom[5125 ] = 12'h8b5;
    rom[5126 ] = 12'h8b5;
    rom[5127 ] = 12'h8b5;
    rom[5128 ] = 12'h8b5;
    rom[5129 ] = 12'h9b5;
    rom[5130 ] = 12'h9b5;
    rom[5131 ] = 12'h9b5;
    rom[5132 ] = 12'h9b5;
    rom[5133 ] = 12'h9b5;
    rom[5134 ] = 12'h9b4;
    rom[5135 ] = 12'h9b4;
    rom[5136 ] = 12'h9b4;
    rom[5137 ] = 12'h9b4;
    rom[5138 ] = 12'h9b4;
    rom[5139 ] = 12'h9b4;
    rom[5140 ] = 12'hab4;
    rom[5141 ] = 12'h000;
    rom[5142 ] = 12'h000;
    rom[5143 ] = 12'h000;
    rom[5144 ] = 12'h000;
    rom[5145 ] = 12'h000;
    rom[5146 ] = 12'h000;
    rom[5147 ] = 12'h000;
    rom[5148 ] = 12'h000;
    rom[5149 ] = 12'h000;
    rom[5150 ] = 12'h000;
    rom[5151 ] = 12'h000;
    rom[5152 ] = 12'h000;
    rom[5153 ] = 12'h000;
    rom[5154 ] = 12'h000;
    rom[5155 ] = 12'h000;
    rom[5156 ] = 12'h000;
    rom[5157 ] = 12'h000;
    rom[5158 ] = 12'h000;
    rom[5159 ] = 12'h000;
    rom[5160 ] = 12'h000;
    rom[5161 ] = 12'h000;
    rom[5162 ] = 12'h000;
    rom[5163 ] = 12'h000;
    rom[5164 ] = 12'h000;
    rom[5165 ] = 12'h000;
    rom[5166 ] = 12'h000;
    rom[5167 ] = 12'h000;
    rom[5168 ] = 12'h000;
    rom[5169 ] = 12'h000;
    rom[5170 ] = 12'h000;
    rom[5171 ] = 12'h000;
    rom[5172 ] = 12'h000;
    rom[5173 ] = 12'h000;
    rom[5174 ] = 12'h000;
    rom[5175 ] = 12'h000;
    rom[5176 ] = 12'h000;
    rom[5177 ] = 12'h000;
    rom[5178 ] = 12'h000;
    rom[5179 ] = 12'h000;
    rom[5180 ] = 12'h000;
    rom[5181 ] = 12'h000;
    rom[5182 ] = 12'h000;
    rom[5183 ] = 12'h000;
    rom[5184 ] = 12'h000;
    rom[5185 ] = 12'h000;
    rom[5186 ] = 12'h000;
    rom[5187 ] = 12'h000;
    rom[5188 ] = 12'h000;
    rom[5189 ] = 12'h000;
    rom[5190 ] = 12'h000;
    rom[5191 ] = 12'h000;
    rom[5192 ] = 12'h000;
    rom[5193 ] = 12'h000;
    rom[5194 ] = 12'h000;
    rom[5195 ] = 12'h000;
    rom[5196 ] = 12'h000;
    rom[5197 ] = 12'h000;
    rom[5198 ] = 12'h000;
    rom[5199 ] = 12'h000;
    rom[5200 ] = 12'h000;
    rom[5201 ] = 12'h000;
    rom[5202 ] = 12'h000;
    rom[5203 ] = 12'h000;
    rom[5204 ] = 12'h000;
    rom[5205 ] = 12'h000;
    rom[5206 ] = 12'h000;
    rom[5207 ] = 12'h000;
    rom[5208 ] = 12'h000;
    rom[5209 ] = 12'h000;
    rom[5210 ] = 12'h000;
    rom[5211 ] = 12'h000;
    rom[5212 ] = 12'h000;
    rom[5213 ] = 12'h3a2;
    rom[5214 ] = 12'h3a2;
    rom[5215 ] = 12'h3a2;
    rom[5216 ] = 12'h3a2;
    rom[5217 ] = 12'h3a2;
    rom[5218 ] = 12'h3a2;
    rom[5219 ] = 12'h3a2;
    rom[5220 ] = 12'h3a2;
    rom[5221 ] = 12'h3a2;
    rom[5222 ] = 12'h3a2;
    rom[5223 ] = 12'h3a2;
    rom[5224 ] = 12'h3a2;
    rom[5225 ] = 12'h3a2;
    rom[5226 ] = 12'h3a2;
    rom[5227 ] = 12'h3a2;
    rom[5228 ] = 12'h3a2;
    rom[5229 ] = 12'h3a2;
    rom[5230 ] = 12'h3a2;
    rom[5231 ] = 12'h3a2;
    rom[5232 ] = 12'h3a2;
    rom[5233 ] = 12'h3a2;
    rom[5234 ] = 12'h3a2;
    rom[5235 ] = 12'h3a2;
    rom[5236 ] = 12'h3a2;
    rom[5237 ] = 12'h3a2;
    rom[5238 ] = 12'h3a2;
    rom[5239 ] = 12'h000;
    rom[5240 ] = 12'h000;
    rom[5241 ] = 12'h000;
    rom[5242 ] = 12'h000;
    rom[5243 ] = 12'h000;
    rom[5244 ] = 12'h000;
    rom[5245 ] = 12'h000;
    rom[5246 ] = 12'h000;
    rom[5247 ] = 12'h000;
    rom[5248 ] = 12'h000;
    rom[5249 ] = 12'h000;
    rom[5250 ] = 12'h000;
    rom[5251 ] = 12'h000;
    rom[5252 ] = 12'h8b6;
    rom[5253 ] = 12'h8b5;
    rom[5254 ] = 12'h8b5;
    rom[5255 ] = 12'h8b5;
    rom[5256 ] = 12'h8b5;
    rom[5257 ] = 12'h8b5;
    rom[5258 ] = 12'h8b5;
    rom[5259 ] = 12'h8b5;
    rom[5260 ] = 12'h9b5;
    rom[5261 ] = 12'h9b5;
    rom[5262 ] = 12'h9b5;
    rom[5263 ] = 12'h9b5;
    rom[5264 ] = 12'h9b5;
    rom[5265 ] = 12'h9b4;
    rom[5266 ] = 12'h9b4;
    rom[5267 ] = 12'h9b4;
    rom[5268 ] = 12'h000;
    rom[5269 ] = 12'h000;
    rom[5270 ] = 12'h000;
    rom[5271 ] = 12'h000;
    rom[5272 ] = 12'h000;
    rom[5273 ] = 12'h000;
    rom[5274 ] = 12'h000;
    rom[5275 ] = 12'h000;
    rom[5276 ] = 12'h000;
    rom[5277 ] = 12'h000;
    rom[5278 ] = 12'h000;
    rom[5279 ] = 12'h000;
    rom[5280 ] = 12'h000;
    rom[5281 ] = 12'h000;
    rom[5282 ] = 12'h000;
    rom[5283 ] = 12'h000;
    rom[5284 ] = 12'h000;
    rom[5285 ] = 12'h000;
    rom[5286 ] = 12'h000;
    rom[5287 ] = 12'h000;
    rom[5288 ] = 12'h000;
    rom[5289 ] = 12'h000;
    rom[5290 ] = 12'h000;
    rom[5291 ] = 12'h000;
    rom[5292 ] = 12'h000;
    rom[5293 ] = 12'h000;
    rom[5294 ] = 12'h000;
    rom[5295 ] = 12'h000;
    rom[5296 ] = 12'h000;
    rom[5297 ] = 12'h000;
    rom[5298 ] = 12'h000;
    rom[5299 ] = 12'h000;
    rom[5300 ] = 12'h000;
    rom[5301 ] = 12'h000;
    rom[5302 ] = 12'h000;
    rom[5303 ] = 12'h000;
    rom[5304 ] = 12'h000;
    rom[5305 ] = 12'h000;
    rom[5306 ] = 12'h000;
    rom[5307 ] = 12'h000;
    rom[5308 ] = 12'h000;
    rom[5309 ] = 12'h000;
    rom[5310 ] = 12'h000;
    rom[5311 ] = 12'h000;
    rom[5312 ] = 12'h000;
    rom[5313 ] = 12'h000;
    rom[5314 ] = 12'h000;
    rom[5315 ] = 12'h000;
    rom[5316 ] = 12'h000;
    rom[5317 ] = 12'h000;
    rom[5318 ] = 12'h000;
    rom[5319 ] = 12'h000;
    rom[5320 ] = 12'h000;
    rom[5321 ] = 12'h000;
    rom[5322 ] = 12'h000;
    rom[5323 ] = 12'h000;
    rom[5324 ] = 12'h000;
    rom[5325 ] = 12'h000;
    rom[5326 ] = 12'h000;
    rom[5327 ] = 12'h000;
    rom[5328 ] = 12'h000;
    rom[5329 ] = 12'h000;
    rom[5330 ] = 12'h000;
    rom[5331 ] = 12'h000;
    rom[5332 ] = 12'h000;
    rom[5333 ] = 12'h000;
    rom[5334 ] = 12'h000;
    rom[5335 ] = 12'h000;
    rom[5336 ] = 12'h000;
    rom[5337 ] = 12'h000;
    rom[5338 ] = 12'h000;
    rom[5339 ] = 12'h000;
    rom[5340 ] = 12'h3a2;
    rom[5341 ] = 12'h3a2;
    rom[5342 ] = 12'h3a2;
    rom[5343 ] = 12'h3a2;
    rom[5344 ] = 12'h3a2;
    rom[5345 ] = 12'h3a2;
    rom[5346 ] = 12'h3a2;
    rom[5347 ] = 12'h3a2;
    rom[5348 ] = 12'h3a2;
    rom[5349 ] = 12'h3a2;
    rom[5350 ] = 12'h3a2;
    rom[5351 ] = 12'h3a2;
    rom[5352 ] = 12'h3a2;
    rom[5353 ] = 12'h3a2;
    rom[5354 ] = 12'h3a2;
    rom[5355 ] = 12'h3a2;
    rom[5356 ] = 12'h3a2;
    rom[5357 ] = 12'h3a2;
    rom[5358 ] = 12'h3a2;
    rom[5359 ] = 12'h3a2;
    rom[5360 ] = 12'h3a2;
    rom[5361 ] = 12'h3a2;
    rom[5362 ] = 12'h3a2;
    rom[5363 ] = 12'h3a2;
    rom[5364 ] = 12'h3a2;
    rom[5365 ] = 12'h000;
    rom[5366 ] = 12'h000;
    rom[5367 ] = 12'h000;
    rom[5368 ] = 12'h000;
    rom[5369 ] = 12'h000;
    rom[5370 ] = 12'h000;
    rom[5371 ] = 12'h000;
    rom[5372 ] = 12'h000;
    rom[5373 ] = 12'h000;
    rom[5374 ] = 12'h000;
    rom[5375 ] = 12'h000;
    rom[5376 ] = 12'h000;
    rom[5377 ] = 12'h000;
    rom[5378 ] = 12'h000;
    rom[5379 ] = 12'h000;
    rom[5380 ] = 12'h8b6;
    rom[5381 ] = 12'h8b6;
    rom[5382 ] = 12'h8b6;
    rom[5383 ] = 12'h8b6;
    rom[5384 ] = 12'h8b5;
    rom[5385 ] = 12'h8b5;
    rom[5386 ] = 12'h8b5;
    rom[5387 ] = 12'h8b5;
    rom[5388 ] = 12'h8b5;
    rom[5389 ] = 12'h8b5;
    rom[5390 ] = 12'h8b5;
    rom[5391 ] = 12'h9b5;
    rom[5392 ] = 12'h9b5;
    rom[5393 ] = 12'h9b5;
    rom[5394 ] = 12'h9b5;
    rom[5395 ] = 12'h9b5;
    rom[5396 ] = 12'h000;
    rom[5397 ] = 12'h000;
    rom[5398 ] = 12'h000;
    rom[5399 ] = 12'h000;
    rom[5400 ] = 12'h000;
    rom[5401 ] = 12'h000;
    rom[5402 ] = 12'h000;
    rom[5403 ] = 12'h000;
    rom[5404 ] = 12'h000;
    rom[5405 ] = 12'h000;
    rom[5406 ] = 12'h000;
    rom[5407 ] = 12'h000;
    rom[5408 ] = 12'h000;
    rom[5409 ] = 12'h000;
    rom[5410 ] = 12'h000;
    rom[5411 ] = 12'h000;
    rom[5412 ] = 12'h000;
    rom[5413 ] = 12'h000;
    rom[5414 ] = 12'h000;
    rom[5415 ] = 12'h000;
    rom[5416 ] = 12'h000;
    rom[5417 ] = 12'h000;
    rom[5418 ] = 12'h000;
    rom[5419 ] = 12'h000;
    rom[5420 ] = 12'h000;
    rom[5421 ] = 12'h000;
    rom[5422 ] = 12'h000;
    rom[5423 ] = 12'h000;
    rom[5424 ] = 12'h000;
    rom[5425 ] = 12'h000;
    rom[5426 ] = 12'h000;
    rom[5427 ] = 12'h000;
    rom[5428 ] = 12'h000;
    rom[5429 ] = 12'h000;
    rom[5430 ] = 12'h000;
    rom[5431 ] = 12'h000;
    rom[5432 ] = 12'h000;
    rom[5433 ] = 12'h000;
    rom[5434 ] = 12'h000;
    rom[5435 ] = 12'h000;
    rom[5436 ] = 12'h000;
    rom[5437 ] = 12'h000;
    rom[5438 ] = 12'h000;
    rom[5439 ] = 12'h000;
    rom[5440 ] = 12'h000;
    rom[5441 ] = 12'h000;
    rom[5442 ] = 12'h000;
    rom[5443 ] = 12'h000;
    rom[5444 ] = 12'h000;
    rom[5445 ] = 12'h000;
    rom[5446 ] = 12'h000;
    rom[5447 ] = 12'h000;
    rom[5448 ] = 12'h000;
    rom[5449 ] = 12'h000;
    rom[5450 ] = 12'h000;
    rom[5451 ] = 12'h000;
    rom[5452 ] = 12'h000;
    rom[5453 ] = 12'h000;
    rom[5454 ] = 12'h000;
    rom[5455 ] = 12'h000;
    rom[5456 ] = 12'h000;
    rom[5457 ] = 12'h000;
    rom[5458 ] = 12'h000;
    rom[5459 ] = 12'h000;
    rom[5460 ] = 12'h000;
    rom[5461 ] = 12'h000;
    rom[5462 ] = 12'h000;
    rom[5463 ] = 12'h000;
    rom[5464 ] = 12'h000;
    rom[5465 ] = 12'h000;
    rom[5466 ] = 12'h000;
    rom[5467 ] = 12'h3a2;
    rom[5468 ] = 12'h3a2;
    rom[5469 ] = 12'h3a2;
    rom[5470 ] = 12'h3a2;
    rom[5471 ] = 12'h3a2;
    rom[5472 ] = 12'h3a2;
    rom[5473 ] = 12'h3a2;
    rom[5474 ] = 12'h3a2;
    rom[5475 ] = 12'h3a2;
    rom[5476 ] = 12'h3a2;
    rom[5477 ] = 12'h3a2;
    rom[5478 ] = 12'h3a2;
    rom[5479 ] = 12'h3a2;
    rom[5480 ] = 12'h3a2;
    rom[5481 ] = 12'h3a2;
    rom[5482 ] = 12'h3a2;
    rom[5483 ] = 12'h3a2;
    rom[5484 ] = 12'h3a2;
    rom[5485 ] = 12'h3a2;
    rom[5486 ] = 12'h3a2;
    rom[5487 ] = 12'h3a2;
    rom[5488 ] = 12'h3a2;
    rom[5489 ] = 12'h3a2;
    rom[5490 ] = 12'h3a2;
    rom[5491 ] = 12'h3a2;
    rom[5492 ] = 12'h000;
    rom[5493 ] = 12'h000;
    rom[5494 ] = 12'h000;
    rom[5495 ] = 12'h000;
    rom[5496 ] = 12'h000;
    rom[5497 ] = 12'h000;
    rom[5498 ] = 12'h000;
    rom[5499 ] = 12'h000;
    rom[5500 ] = 12'h000;
    rom[5501 ] = 12'h000;
    rom[5502 ] = 12'h000;
    rom[5503 ] = 12'h000;
    rom[5504 ] = 12'h000;
    rom[5505 ] = 12'h000;
    rom[5506 ] = 12'h000;
    rom[5507 ] = 12'h7b6;
    rom[5508 ] = 12'h7b6;
    rom[5509 ] = 12'h7b6;
    rom[5510 ] = 12'h7b6;
    rom[5511 ] = 12'h8b6;
    rom[5512 ] = 12'h8b6;
    rom[5513 ] = 12'h8b6;
    rom[5514 ] = 12'h8b5;
    rom[5515 ] = 12'h8b5;
    rom[5516 ] = 12'h8b5;
    rom[5517 ] = 12'h8b5;
    rom[5518 ] = 12'h8b5;
    rom[5519 ] = 12'h8b5;
    rom[5520 ] = 12'h8b5;
    rom[5521 ] = 12'h9b5;
    rom[5522 ] = 12'h9b5;
    rom[5523 ] = 12'h000;
    rom[5524 ] = 12'h000;
    rom[5525 ] = 12'h000;
    rom[5526 ] = 12'h000;
    rom[5527 ] = 12'h000;
    rom[5528 ] = 12'h000;
    rom[5529 ] = 12'h000;
    rom[5530 ] = 12'h000;
    rom[5531 ] = 12'h000;
    rom[5532 ] = 12'h000;
    rom[5533 ] = 12'h000;
    rom[5534 ] = 12'h000;
    rom[5535 ] = 12'h000;
    rom[5536 ] = 12'h000;
    rom[5537 ] = 12'h000;
    rom[5538 ] = 12'h000;
    rom[5539 ] = 12'h000;
    rom[5540 ] = 12'h000;
    rom[5541 ] = 12'h000;
    rom[5542 ] = 12'h000;
    rom[5543 ] = 12'h000;
    rom[5544 ] = 12'h000;
    rom[5545 ] = 12'h000;
    rom[5546 ] = 12'h000;
    rom[5547 ] = 12'h000;
    rom[5548 ] = 12'h000;
    rom[5549 ] = 12'h000;
    rom[5550 ] = 12'h000;
    rom[5551 ] = 12'h000;
    rom[5552 ] = 12'h000;
    rom[5553 ] = 12'h000;
    rom[5554 ] = 12'h000;
    rom[5555 ] = 12'h000;
    rom[5556 ] = 12'h000;
    rom[5557 ] = 12'h000;
    rom[5558 ] = 12'h000;
    rom[5559 ] = 12'h000;
    rom[5560 ] = 12'h000;
    rom[5561 ] = 12'h000;
    rom[5562 ] = 12'h000;
    rom[5563 ] = 12'h000;
    rom[5564 ] = 12'h000;
    rom[5565 ] = 12'h000;
    rom[5566 ] = 12'h000;
    rom[5567 ] = 12'h000;
    rom[5568 ] = 12'h000;
    rom[5569 ] = 12'h000;
    rom[5570 ] = 12'h000;
    rom[5571 ] = 12'h000;
    rom[5572 ] = 12'h000;
    rom[5573 ] = 12'h000;
    rom[5574 ] = 12'h000;
    rom[5575 ] = 12'h000;
    rom[5576 ] = 12'h000;
    rom[5577 ] = 12'h000;
    rom[5578 ] = 12'h000;
    rom[5579 ] = 12'h000;
    rom[5580 ] = 12'h000;
    rom[5581 ] = 12'h000;
    rom[5582 ] = 12'h000;
    rom[5583 ] = 12'h000;
    rom[5584 ] = 12'h000;
    rom[5585 ] = 12'h000;
    rom[5586 ] = 12'h000;
    rom[5587 ] = 12'h000;
    rom[5588 ] = 12'h000;
    rom[5589 ] = 12'h000;
    rom[5590 ] = 12'h000;
    rom[5591 ] = 12'h000;
    rom[5592 ] = 12'h000;
    rom[5593 ] = 12'h3a2;
    rom[5594 ] = 12'h3a2;
    rom[5595 ] = 12'h3a2;
    rom[5596 ] = 12'h3a2;
    rom[5597 ] = 12'h3a2;
    rom[5598 ] = 12'h3a2;
    rom[5599 ] = 12'h3a2;
    rom[5600 ] = 12'h3a2;
    rom[5601 ] = 12'h3a2;
    rom[5602 ] = 12'h3a2;
    rom[5603 ] = 12'h3a2;
    rom[5604 ] = 12'h3a2;
    rom[5605 ] = 12'h3a2;
    rom[5606 ] = 12'h3a2;
    rom[5607 ] = 12'h3a2;
    rom[5608 ] = 12'h3a2;
    rom[5609 ] = 12'h3a2;
    rom[5610 ] = 12'h3a2;
    rom[5611 ] = 12'h3a2;
    rom[5612 ] = 12'h3a2;
    rom[5613 ] = 12'h3a2;
    rom[5614 ] = 12'h3a2;
    rom[5615 ] = 12'h3a2;
    rom[5616 ] = 12'h3a2;
    rom[5617 ] = 12'h3a2;
    rom[5618 ] = 12'h392;
    rom[5619 ] = 12'h000;
    rom[5620 ] = 12'h000;
    rom[5621 ] = 12'h000;
    rom[5622 ] = 12'h000;
    rom[5623 ] = 12'h000;
    rom[5624 ] = 12'h000;
    rom[5625 ] = 12'h000;
    rom[5626 ] = 12'h000;
    rom[5627 ] = 12'h000;
    rom[5628 ] = 12'h000;
    rom[5629 ] = 12'h000;
    rom[5630 ] = 12'h000;
    rom[5631 ] = 12'h000;
    rom[5632 ] = 12'h000;
    rom[5633 ] = 12'h000;
    rom[5634 ] = 12'h000;
    rom[5635 ] = 12'h7c6;
    rom[5636 ] = 12'h7b6;
    rom[5637 ] = 12'h7b6;
    rom[5638 ] = 12'h7b6;
    rom[5639 ] = 12'h7b6;
    rom[5640 ] = 12'h7b6;
    rom[5641 ] = 12'h7b6;
    rom[5642 ] = 12'h8b6;
    rom[5643 ] = 12'h8b6;
    rom[5644 ] = 12'h8b6;
    rom[5645 ] = 12'h8b5;
    rom[5646 ] = 12'h8b5;
    rom[5647 ] = 12'h8b5;
    rom[5648 ] = 12'h8b5;
    rom[5649 ] = 12'h8b5;
    rom[5650 ] = 12'h8b5;
    rom[5651 ] = 12'h000;
    rom[5652 ] = 12'h000;
    rom[5653 ] = 12'h000;
    rom[5654 ] = 12'h000;
    rom[5655 ] = 12'h000;
    rom[5656 ] = 12'h000;
    rom[5657 ] = 12'h000;
    rom[5658 ] = 12'h000;
    rom[5659 ] = 12'h000;
    rom[5660 ] = 12'h000;
    rom[5661 ] = 12'h000;
    rom[5662 ] = 12'h000;
    rom[5663 ] = 12'h000;
    rom[5664 ] = 12'h000;
    rom[5665 ] = 12'h000;
    rom[5666 ] = 12'h000;
    rom[5667 ] = 12'h000;
    rom[5668 ] = 12'h000;
    rom[5669 ] = 12'h000;
    rom[5670 ] = 12'h000;
    rom[5671 ] = 12'h000;
    rom[5672 ] = 12'h000;
    rom[5673 ] = 12'h000;
    rom[5674 ] = 12'h000;
    rom[5675 ] = 12'h000;
    rom[5676 ] = 12'h000;
    rom[5677 ] = 12'h000;
    rom[5678 ] = 12'h000;
    rom[5679 ] = 12'h000;
    rom[5680 ] = 12'h000;
    rom[5681 ] = 12'h000;
    rom[5682 ] = 12'h000;
    rom[5683 ] = 12'h000;
    rom[5684 ] = 12'h000;
    rom[5685 ] = 12'h000;
    rom[5686 ] = 12'h000;
    rom[5687 ] = 12'h000;
    rom[5688 ] = 12'h000;
    rom[5689 ] = 12'h000;
    rom[5690 ] = 12'h000;
    rom[5691 ] = 12'h000;
    rom[5692 ] = 12'h000;
    rom[5693 ] = 12'h000;
    rom[5694 ] = 12'h000;
    rom[5695 ] = 12'h000;
    rom[5696 ] = 12'h000;
    rom[5697 ] = 12'h000;
    rom[5698 ] = 12'h000;
    rom[5699 ] = 12'h000;
    rom[5700 ] = 12'h000;
    rom[5701 ] = 12'h000;
    rom[5702 ] = 12'h000;
    rom[5703 ] = 12'h000;
    rom[5704 ] = 12'h000;
    rom[5705 ] = 12'h000;
    rom[5706 ] = 12'h000;
    rom[5707 ] = 12'h000;
    rom[5708 ] = 12'h000;
    rom[5709 ] = 12'h000;
    rom[5710 ] = 12'h000;
    rom[5711 ] = 12'h000;
    rom[5712 ] = 12'h000;
    rom[5713 ] = 12'h000;
    rom[5714 ] = 12'h000;
    rom[5715 ] = 12'h000;
    rom[5716 ] = 12'h000;
    rom[5717 ] = 12'h000;
    rom[5718 ] = 12'h000;
    rom[5719 ] = 12'h000;
    rom[5720 ] = 12'h3a2;
    rom[5721 ] = 12'h3a2;
    rom[5722 ] = 12'h3a2;
    rom[5723 ] = 12'h3a2;
    rom[5724 ] = 12'h3a2;
    rom[5725 ] = 12'h3a2;
    rom[5726 ] = 12'h3a2;
    rom[5727 ] = 12'h3a2;
    rom[5728 ] = 12'h3a2;
    rom[5729 ] = 12'h3a2;
    rom[5730 ] = 12'h3a2;
    rom[5731 ] = 12'h3a2;
    rom[5732 ] = 12'h3a2;
    rom[5733 ] = 12'h3a2;
    rom[5734 ] = 12'h3a2;
    rom[5735 ] = 12'h3a2;
    rom[5736 ] = 12'h3a2;
    rom[5737 ] = 12'h3a2;
    rom[5738 ] = 12'h3a2;
    rom[5739 ] = 12'h3a2;
    rom[5740 ] = 12'h3a2;
    rom[5741 ] = 12'h3a2;
    rom[5742 ] = 12'h3a2;
    rom[5743 ] = 12'h3a2;
    rom[5744 ] = 12'h3a2;
    rom[5745 ] = 12'h000;
    rom[5746 ] = 12'h000;
    rom[5747 ] = 12'h000;
    rom[5748 ] = 12'h000;
    rom[5749 ] = 12'h000;
    rom[5750 ] = 12'h000;
    rom[5751 ] = 12'h000;
    rom[5752 ] = 12'h000;
    rom[5753 ] = 12'h000;
    rom[5754 ] = 12'h000;
    rom[5755 ] = 12'h000;
    rom[5756 ] = 12'h000;
    rom[5757 ] = 12'h000;
    rom[5758 ] = 12'h000;
    rom[5759 ] = 12'h000;
    rom[5760 ] = 12'h000;
    rom[5761 ] = 12'h000;
    rom[5762 ] = 12'h000;
    rom[5763 ] = 12'h7c7;
    rom[5764 ] = 12'h7c6;
    rom[5765 ] = 12'h7c6;
    rom[5766 ] = 12'h7c6;
    rom[5767 ] = 12'h7b6;
    rom[5768 ] = 12'h7b6;
    rom[5769 ] = 12'h7b6;
    rom[5770 ] = 12'h7b6;
    rom[5771 ] = 12'h7b6;
    rom[5772 ] = 12'h8b6;
    rom[5773 ] = 12'h8b6;
    rom[5774 ] = 12'h8b6;
    rom[5775 ] = 12'h8b6;
    rom[5776 ] = 12'h8b5;
    rom[5777 ] = 12'h8b5;
    rom[5778 ] = 12'h8b5;
    rom[5779 ] = 12'h000;
    rom[5780 ] = 12'h000;
    rom[5781 ] = 12'h000;
    rom[5782 ] = 12'h000;
    rom[5783 ] = 12'h000;
    rom[5784 ] = 12'h000;
    rom[5785 ] = 12'h000;
    rom[5786 ] = 12'h000;
    rom[5787 ] = 12'h000;
    rom[5788 ] = 12'h000;
    rom[5789 ] = 12'h000;
    rom[5790 ] = 12'h000;
    rom[5791 ] = 12'h000;
    rom[5792 ] = 12'h000;
    rom[5793 ] = 12'h000;
    rom[5794 ] = 12'h000;
    rom[5795 ] = 12'h000;
    rom[5796 ] = 12'h000;
    rom[5797 ] = 12'h000;
    rom[5798 ] = 12'h000;
    rom[5799 ] = 12'h000;
    rom[5800 ] = 12'h000;
    rom[5801 ] = 12'h000;
    rom[5802 ] = 12'h000;
    rom[5803 ] = 12'h000;
    rom[5804 ] = 12'h000;
    rom[5805 ] = 12'h000;
    rom[5806 ] = 12'h000;
    rom[5807 ] = 12'h000;
    rom[5808 ] = 12'h000;
    rom[5809 ] = 12'h000;
    rom[5810 ] = 12'h000;
    rom[5811 ] = 12'h000;
    rom[5812 ] = 12'h000;
    rom[5813 ] = 12'h000;
    rom[5814 ] = 12'h000;
    rom[5815 ] = 12'h000;
    rom[5816 ] = 12'h000;
    rom[5817 ] = 12'h000;
    rom[5818 ] = 12'h000;
    rom[5819 ] = 12'h000;
    rom[5820 ] = 12'h000;
    rom[5821 ] = 12'h000;
    rom[5822 ] = 12'h000;
    rom[5823 ] = 12'h000;
    rom[5824 ] = 12'h000;
    rom[5825 ] = 12'h000;
    rom[5826 ] = 12'h000;
    rom[5827 ] = 12'h000;
    rom[5828 ] = 12'h000;
    rom[5829 ] = 12'h000;
    rom[5830 ] = 12'h000;
    rom[5831 ] = 12'h000;
    rom[5832 ] = 12'h000;
    rom[5833 ] = 12'h000;
    rom[5834 ] = 12'h000;
    rom[5835 ] = 12'h000;
    rom[5836 ] = 12'h000;
    rom[5837 ] = 12'h000;
    rom[5838 ] = 12'h000;
    rom[5839 ] = 12'h000;
    rom[5840 ] = 12'h000;
    rom[5841 ] = 12'h000;
    rom[5842 ] = 12'h000;
    rom[5843 ] = 12'h000;
    rom[5844 ] = 12'h000;
    rom[5845 ] = 12'h000;
    rom[5846 ] = 12'h492;
    rom[5847 ] = 12'h3a2;
    rom[5848 ] = 12'h3a2;
    rom[5849 ] = 12'h3a2;
    rom[5850 ] = 12'h3a2;
    rom[5851 ] = 12'h3a2;
    rom[5852 ] = 12'h3a2;
    rom[5853 ] = 12'h3a2;
    rom[5854 ] = 12'h3a2;
    rom[5855 ] = 12'h3a2;
    rom[5856 ] = 12'h3a2;
    rom[5857 ] = 12'h3a2;
    rom[5858 ] = 12'h3a2;
    rom[5859 ] = 12'h3a2;
    rom[5860 ] = 12'h3a2;
    rom[5861 ] = 12'h3a2;
    rom[5862 ] = 12'h3a2;
    rom[5863 ] = 12'h3a2;
    rom[5864 ] = 12'h3a2;
    rom[5865 ] = 12'h3a2;
    rom[5866 ] = 12'h3a2;
    rom[5867 ] = 12'h3a2;
    rom[5868 ] = 12'h3a2;
    rom[5869 ] = 12'h3a2;
    rom[5870 ] = 12'h3a2;
    rom[5871 ] = 12'h3a2;
    rom[5872 ] = 12'h000;
    rom[5873 ] = 12'h000;
    rom[5874 ] = 12'h000;
    rom[5875 ] = 12'h000;
    rom[5876 ] = 12'h000;
    rom[5877 ] = 12'h000;
    rom[5878 ] = 12'h000;
    rom[5879 ] = 12'h000;
    rom[5880 ] = 12'h000;
    rom[5881 ] = 12'h000;
    rom[5882 ] = 12'h000;
    rom[5883 ] = 12'h000;
    rom[5884 ] = 12'h000;
    rom[5885 ] = 12'h000;
    rom[5886 ] = 12'h000;
    rom[5887 ] = 12'h000;
    rom[5888 ] = 12'h000;
    rom[5889 ] = 12'h000;
    rom[5890 ] = 12'h6c7;
    rom[5891 ] = 12'h6c7;
    rom[5892 ] = 12'h7c7;
    rom[5893 ] = 12'h7c7;
    rom[5894 ] = 12'h7c6;
    rom[5895 ] = 12'h7c6;
    rom[5896 ] = 12'h7c6;
    rom[5897 ] = 12'h7b6;
    rom[5898 ] = 12'h7b6;
    rom[5899 ] = 12'h7b6;
    rom[5900 ] = 12'h7b6;
    rom[5901 ] = 12'h7b6;
    rom[5902 ] = 12'h7b6;
    rom[5903 ] = 12'h8b6;
    rom[5904 ] = 12'h8b6;
    rom[5905 ] = 12'h8b6;
    rom[5906 ] = 12'h000;
    rom[5907 ] = 12'h000;
    rom[5908 ] = 12'h000;
    rom[5909 ] = 12'h000;
    rom[5910 ] = 12'h000;
    rom[5911 ] = 12'h000;
    rom[5912 ] = 12'h000;
    rom[5913 ] = 12'h000;
    rom[5914 ] = 12'h000;
    rom[5915 ] = 12'h000;
    rom[5916 ] = 12'h000;
    rom[5917 ] = 12'h000;
    rom[5918 ] = 12'h000;
    rom[5919 ] = 12'h000;
    rom[5920 ] = 12'h000;
    rom[5921 ] = 12'h000;
    rom[5922 ] = 12'h000;
    rom[5923 ] = 12'h000;
    rom[5924 ] = 12'h000;
    rom[5925 ] = 12'h000;
    rom[5926 ] = 12'h000;
    rom[5927 ] = 12'h000;
    rom[5928 ] = 12'h000;
    rom[5929 ] = 12'h000;
    rom[5930 ] = 12'h000;
    rom[5931 ] = 12'h000;
    rom[5932 ] = 12'h000;
    rom[5933 ] = 12'h000;
    rom[5934 ] = 12'h000;
    rom[5935 ] = 12'h000;
    rom[5936 ] = 12'h000;
    rom[5937 ] = 12'h000;
    rom[5938 ] = 12'h000;
    rom[5939 ] = 12'h000;
    rom[5940 ] = 12'h000;
    rom[5941 ] = 12'h000;
    rom[5942 ] = 12'h000;
    rom[5943 ] = 12'h000;
    rom[5944 ] = 12'h000;
    rom[5945 ] = 12'h000;
    rom[5946 ] = 12'h000;
    rom[5947 ] = 12'h000;
    rom[5948 ] = 12'h000;
    rom[5949 ] = 12'h000;
    rom[5950 ] = 12'h000;
    rom[5951 ] = 12'h000;
    rom[5952 ] = 12'h000;
    rom[5953 ] = 12'h000;
    rom[5954 ] = 12'h000;
    rom[5955 ] = 12'h000;
    rom[5956 ] = 12'h000;
    rom[5957 ] = 12'h000;
    rom[5958 ] = 12'h000;
    rom[5959 ] = 12'h000;
    rom[5960 ] = 12'h000;
    rom[5961 ] = 12'h000;
    rom[5962 ] = 12'h000;
    rom[5963 ] = 12'h000;
    rom[5964 ] = 12'h000;
    rom[5965 ] = 12'h000;
    rom[5966 ] = 12'h000;
    rom[5967 ] = 12'h000;
    rom[5968 ] = 12'h000;
    rom[5969 ] = 12'h000;
    rom[5970 ] = 12'h000;
    rom[5971 ] = 12'h000;
    rom[5972 ] = 12'h000;
    rom[5973 ] = 12'h3a2;
    rom[5974 ] = 12'h3a2;
    rom[5975 ] = 12'h3a2;
    rom[5976 ] = 12'h3a2;
    rom[5977 ] = 12'h3a2;
    rom[5978 ] = 12'h3a2;
    rom[5979 ] = 12'h3a2;
    rom[5980 ] = 12'h3a2;
    rom[5981 ] = 12'h3a2;
    rom[5982 ] = 12'h3a2;
    rom[5983 ] = 12'h3a2;
    rom[5984 ] = 12'h3a2;
    rom[5985 ] = 12'h3a2;
    rom[5986 ] = 12'h3a2;
    rom[5987 ] = 12'h3a2;
    rom[5988 ] = 12'h3a2;
    rom[5989 ] = 12'h3a2;
    rom[5990 ] = 12'h3a2;
    rom[5991 ] = 12'h3a2;
    rom[5992 ] = 12'h3a2;
    rom[5993 ] = 12'h3a2;
    rom[5994 ] = 12'h3a2;
    rom[5995 ] = 12'h3a2;
    rom[5996 ] = 12'h3a2;
    rom[5997 ] = 12'h3a2;
    rom[5998 ] = 12'h4a1;
    rom[5999 ] = 12'h000;
    rom[6000 ] = 12'h000;
    rom[6001 ] = 12'h000;
    rom[6002 ] = 12'h000;
    rom[6003 ] = 12'h000;
    rom[6004 ] = 12'h000;
    rom[6005 ] = 12'h000;
    rom[6006 ] = 12'h000;
    rom[6007 ] = 12'h000;
    rom[6008 ] = 12'h000;
    rom[6009 ] = 12'h000;
    rom[6010 ] = 12'h000;
    rom[6011 ] = 12'h000;
    rom[6012 ] = 12'h000;
    rom[6013 ] = 12'h000;
    rom[6014 ] = 12'h000;
    rom[6015 ] = 12'h000;
    rom[6016 ] = 12'h000;
    rom[6017 ] = 12'h000;
    rom[6018 ] = 12'h6c7;
    rom[6019 ] = 12'h6c7;
    rom[6020 ] = 12'h6c7;
    rom[6021 ] = 12'h6c7;
    rom[6022 ] = 12'h6c7;
    rom[6023 ] = 12'h7c7;
    rom[6024 ] = 12'h7c7;
    rom[6025 ] = 12'h7c6;
    rom[6026 ] = 12'h7c6;
    rom[6027 ] = 12'h7c6;
    rom[6028 ] = 12'h7b6;
    rom[6029 ] = 12'h7b6;
    rom[6030 ] = 12'h7b6;
    rom[6031 ] = 12'h7b6;
    rom[6032 ] = 12'h7b6;
    rom[6033 ] = 12'h8b6;
    rom[6034 ] = 12'h000;
    rom[6035 ] = 12'h000;
    rom[6036 ] = 12'h000;
    rom[6037 ] = 12'h000;
    rom[6038 ] = 12'h000;
    rom[6039 ] = 12'h000;
    rom[6040 ] = 12'h000;
    rom[6041 ] = 12'h000;
    rom[6042 ] = 12'h000;
    rom[6043 ] = 12'h000;
    rom[6044 ] = 12'h000;
    rom[6045 ] = 12'h000;
    rom[6046 ] = 12'h000;
    rom[6047 ] = 12'h000;
    rom[6048 ] = 12'h000;
    rom[6049 ] = 12'h000;
    rom[6050 ] = 12'h000;
    rom[6051 ] = 12'h000;
    rom[6052 ] = 12'h000;
    rom[6053 ] = 12'h000;
    rom[6054 ] = 12'h000;
    rom[6055 ] = 12'h492;
    rom[6056 ] = 12'h3a2;
    rom[6057 ] = 12'h000;
    rom[6058 ] = 12'h000;
    rom[6059 ] = 12'h000;
    rom[6060 ] = 12'h000;
    rom[6061 ] = 12'h000;
    rom[6062 ] = 12'h000;
    rom[6063 ] = 12'h000;
    rom[6064 ] = 12'h000;
    rom[6065 ] = 12'h000;
    rom[6066 ] = 12'h000;
    rom[6067 ] = 12'h000;
    rom[6068 ] = 12'h000;
    rom[6069 ] = 12'h000;
    rom[6070 ] = 12'h000;
    rom[6071 ] = 12'h000;
    rom[6072 ] = 12'h000;
    rom[6073 ] = 12'h000;
    rom[6074 ] = 12'h000;
    rom[6075 ] = 12'h000;
    rom[6076 ] = 12'h000;
    rom[6077 ] = 12'h000;
    rom[6078 ] = 12'h000;
    rom[6079 ] = 12'h000;
    rom[6080 ] = 12'h000;
    rom[6081 ] = 12'h000;
    rom[6082 ] = 12'h000;
    rom[6083 ] = 12'h000;
    rom[6084 ] = 12'h000;
    rom[6085 ] = 12'h000;
    rom[6086 ] = 12'h000;
    rom[6087 ] = 12'h000;
    rom[6088 ] = 12'h000;
    rom[6089 ] = 12'h000;
    rom[6090 ] = 12'h000;
    rom[6091 ] = 12'h000;
    rom[6092 ] = 12'h000;
    rom[6093 ] = 12'h000;
    rom[6094 ] = 12'h000;
    rom[6095 ] = 12'h000;
    rom[6096 ] = 12'h000;
    rom[6097 ] = 12'h000;
    rom[6098 ] = 12'h000;
    rom[6099 ] = 12'h000;
    rom[6100 ] = 12'h3a2;
    rom[6101 ] = 12'h3a2;
    rom[6102 ] = 12'h3a2;
    rom[6103 ] = 12'h3a2;
    rom[6104 ] = 12'h3a2;
    rom[6105 ] = 12'h3a2;
    rom[6106 ] = 12'h3a2;
    rom[6107 ] = 12'h3a2;
    rom[6108 ] = 12'h3a2;
    rom[6109 ] = 12'h3a2;
    rom[6110 ] = 12'h3a2;
    rom[6111 ] = 12'h3a2;
    rom[6112 ] = 12'h3a2;
    rom[6113 ] = 12'h3a2;
    rom[6114 ] = 12'h3a2;
    rom[6115 ] = 12'h3a2;
    rom[6116 ] = 12'h3a2;
    rom[6117 ] = 12'h3a2;
    rom[6118 ] = 12'h3a2;
    rom[6119 ] = 12'h3a2;
    rom[6120 ] = 12'h3a2;
    rom[6121 ] = 12'h3a2;
    rom[6122 ] = 12'h3a2;
    rom[6123 ] = 12'h3a2;
    rom[6124 ] = 12'h3a2;
    rom[6125 ] = 12'h000;
    rom[6126 ] = 12'h000;
    rom[6127 ] = 12'h000;
    rom[6128 ] = 12'h000;
    rom[6129 ] = 12'h000;
    rom[6130 ] = 12'h000;
    rom[6131 ] = 12'h000;
    rom[6132 ] = 12'h000;
    rom[6133 ] = 12'h000;
    rom[6134 ] = 12'h000;
    rom[6135 ] = 12'h000;
    rom[6136 ] = 12'h000;
    rom[6137 ] = 12'h000;
    rom[6138 ] = 12'h000;
    rom[6139 ] = 12'h000;
    rom[6140 ] = 12'h000;
    rom[6141 ] = 12'h000;
    rom[6142 ] = 12'h000;
    rom[6143 ] = 12'h000;
    rom[6144 ] = 12'h000;
    rom[6145 ] = 12'h000;
    rom[6146 ] = 12'h6c7;
    rom[6147 ] = 12'h6c7;
    rom[6148 ] = 12'h6c7;
    rom[6149 ] = 12'h6c7;
    rom[6150 ] = 12'h6c7;
    rom[6151 ] = 12'h6c7;
    rom[6152 ] = 12'h6c7;
    rom[6153 ] = 12'h7c7;
    rom[6154 ] = 12'h7c7;
    rom[6155 ] = 12'h7c7;
    rom[6156 ] = 12'h7c6;
    rom[6157 ] = 12'h7c6;
    rom[6158 ] = 12'h7c6;
    rom[6159 ] = 12'h7b6;
    rom[6160 ] = 12'h7b6;
    rom[6161 ] = 12'h000;
    rom[6162 ] = 12'h000;
    rom[6163 ] = 12'h000;
    rom[6164 ] = 12'h000;
    rom[6165 ] = 12'h000;
    rom[6166 ] = 12'h000;
    rom[6167 ] = 12'h000;
    rom[6168 ] = 12'h000;
    rom[6169 ] = 12'h000;
    rom[6170 ] = 12'h000;
    rom[6171 ] = 12'h000;
    rom[6172 ] = 12'h000;
    rom[6173 ] = 12'h000;
    rom[6174 ] = 12'h000;
    rom[6175 ] = 12'h000;
    rom[6176 ] = 12'h000;
    rom[6177 ] = 12'h000;
    rom[6178 ] = 12'h000;
    rom[6179 ] = 12'h000;
    rom[6180 ] = 12'h000;
    rom[6181 ] = 12'h000;
    rom[6182 ] = 12'h000;
    rom[6183 ] = 12'h492;
    rom[6184 ] = 12'h3a2;
    rom[6185 ] = 12'h3a2;
    rom[6186 ] = 12'h000;
    rom[6187 ] = 12'h000;
    rom[6188 ] = 12'h000;
    rom[6189 ] = 12'h000;
    rom[6190 ] = 12'h000;
    rom[6191 ] = 12'h000;
    rom[6192 ] = 12'h000;
    rom[6193 ] = 12'h000;
    rom[6194 ] = 12'h000;
    rom[6195 ] = 12'h000;
    rom[6196 ] = 12'h000;
    rom[6197 ] = 12'h000;
    rom[6198 ] = 12'h000;
    rom[6199 ] = 12'h000;
    rom[6200 ] = 12'h000;
    rom[6201 ] = 12'h000;
    rom[6202 ] = 12'h000;
    rom[6203 ] = 12'h000;
    rom[6204 ] = 12'h000;
    rom[6205 ] = 12'h000;
    rom[6206 ] = 12'h000;
    rom[6207 ] = 12'h000;
    rom[6208 ] = 12'h000;
    rom[6209 ] = 12'h000;
    rom[6210 ] = 12'h000;
    rom[6211 ] = 12'h000;
    rom[6212 ] = 12'h000;
    rom[6213 ] = 12'h000;
    rom[6214 ] = 12'h000;
    rom[6215 ] = 12'h000;
    rom[6216 ] = 12'h000;
    rom[6217 ] = 12'h000;
    rom[6218 ] = 12'h000;
    rom[6219 ] = 12'h000;
    rom[6220 ] = 12'h000;
    rom[6221 ] = 12'h000;
    rom[6222 ] = 12'h000;
    rom[6223 ] = 12'h000;
    rom[6224 ] = 12'h000;
    rom[6225 ] = 12'h000;
    rom[6226 ] = 12'h3a2;
    rom[6227 ] = 12'h3a2;
    rom[6228 ] = 12'h3a2;
    rom[6229 ] = 12'h3a2;
    rom[6230 ] = 12'h3a2;
    rom[6231 ] = 12'h3a2;
    rom[6232 ] = 12'h3a2;
    rom[6233 ] = 12'h3a2;
    rom[6234 ] = 12'h3a2;
    rom[6235 ] = 12'h3a2;
    rom[6236 ] = 12'h3a2;
    rom[6237 ] = 12'h3a2;
    rom[6238 ] = 12'h3a2;
    rom[6239 ] = 12'h3a2;
    rom[6240 ] = 12'h3a2;
    rom[6241 ] = 12'h3a2;
    rom[6242 ] = 12'h3a2;
    rom[6243 ] = 12'h3a2;
    rom[6244 ] = 12'h3a2;
    rom[6245 ] = 12'h3a2;
    rom[6246 ] = 12'h3a2;
    rom[6247 ] = 12'h3a2;
    rom[6248 ] = 12'h3a2;
    rom[6249 ] = 12'h3a2;
    rom[6250 ] = 12'h3a2;
    rom[6251 ] = 12'h3a2;
    rom[6252 ] = 12'h000;
    rom[6253 ] = 12'h000;
    rom[6254 ] = 12'h000;
    rom[6255 ] = 12'h000;
    rom[6256 ] = 12'h000;
    rom[6257 ] = 12'h000;
    rom[6258 ] = 12'h000;
    rom[6259 ] = 12'h000;
    rom[6260 ] = 12'h000;
    rom[6261 ] = 12'h000;
    rom[6262 ] = 12'h000;
    rom[6263 ] = 12'h000;
    rom[6264 ] = 12'h000;
    rom[6265 ] = 12'h000;
    rom[6266 ] = 12'h000;
    rom[6267 ] = 12'h000;
    rom[6268 ] = 12'h000;
    rom[6269 ] = 12'h000;
    rom[6270 ] = 12'h000;
    rom[6271 ] = 12'h000;
    rom[6272 ] = 12'h000;
    rom[6273 ] = 12'h000;
    rom[6274 ] = 12'h6c8;
    rom[6275 ] = 12'h6c7;
    rom[6276 ] = 12'h6c7;
    rom[6277 ] = 12'h6c7;
    rom[6278 ] = 12'h6c7;
    rom[6279 ] = 12'h6c7;
    rom[6280 ] = 12'h6c7;
    rom[6281 ] = 12'h6c7;
    rom[6282 ] = 12'h6c7;
    rom[6283 ] = 12'h6c7;
    rom[6284 ] = 12'h7c7;
    rom[6285 ] = 12'h7c7;
    rom[6286 ] = 12'h7c6;
    rom[6287 ] = 12'h7c6;
    rom[6288 ] = 12'h7c6;
    rom[6289 ] = 12'h000;
    rom[6290 ] = 12'h000;
    rom[6291 ] = 12'h000;
    rom[6292 ] = 12'h000;
    rom[6293 ] = 12'h000;
    rom[6294 ] = 12'h000;
    rom[6295 ] = 12'h000;
    rom[6296 ] = 12'h000;
    rom[6297 ] = 12'h000;
    rom[6298 ] = 12'h000;
    rom[6299 ] = 12'h000;
    rom[6300 ] = 12'h000;
    rom[6301 ] = 12'h000;
    rom[6302 ] = 12'h000;
    rom[6303 ] = 12'h000;
    rom[6304 ] = 12'h000;
    rom[6305 ] = 12'h000;
    rom[6306 ] = 12'h000;
    rom[6307 ] = 12'h000;
    rom[6308 ] = 12'h000;
    rom[6309 ] = 12'h000;
    rom[6310 ] = 12'h000;
    rom[6311 ] = 12'h492;
    rom[6312 ] = 12'h3a2;
    rom[6313 ] = 12'h3a2;
    rom[6314 ] = 12'h3a2;
    rom[6315 ] = 12'h3a2;
    rom[6316 ] = 12'h000;
    rom[6317 ] = 12'h000;
    rom[6318 ] = 12'h000;
    rom[6319 ] = 12'h000;
    rom[6320 ] = 12'h000;
    rom[6321 ] = 12'h000;
    rom[6322 ] = 12'h000;
    rom[6323 ] = 12'h000;
    rom[6324 ] = 12'h000;
    rom[6325 ] = 12'h000;
    rom[6326 ] = 12'h000;
    rom[6327 ] = 12'h000;
    rom[6328 ] = 12'h000;
    rom[6329 ] = 12'h000;
    rom[6330 ] = 12'h000;
    rom[6331 ] = 12'h000;
    rom[6332 ] = 12'h000;
    rom[6333 ] = 12'h000;
    rom[6334 ] = 12'h000;
    rom[6335 ] = 12'h000;
    rom[6336 ] = 12'h000;
    rom[6337 ] = 12'h000;
    rom[6338 ] = 12'h000;
    rom[6339 ] = 12'h000;
    rom[6340 ] = 12'h000;
    rom[6341 ] = 12'h000;
    rom[6342 ] = 12'h000;
    rom[6343 ] = 12'h000;
    rom[6344 ] = 12'h000;
    rom[6345 ] = 12'h000;
    rom[6346 ] = 12'h000;
    rom[6347 ] = 12'h000;
    rom[6348 ] = 12'h000;
    rom[6349 ] = 12'h000;
    rom[6350 ] = 12'h000;
    rom[6351 ] = 12'h000;
    rom[6352 ] = 12'h000;
    rom[6353 ] = 12'h3a2;
    rom[6354 ] = 12'h3a2;
    rom[6355 ] = 12'h3a2;
    rom[6356 ] = 12'h3a2;
    rom[6357 ] = 12'h3a2;
    rom[6358 ] = 12'h3a2;
    rom[6359 ] = 12'h3a2;
    rom[6360 ] = 12'h3a2;
    rom[6361 ] = 12'h3a2;
    rom[6362 ] = 12'h3a2;
    rom[6363 ] = 12'h3a2;
    rom[6364 ] = 12'h3a2;
    rom[6365 ] = 12'h3a2;
    rom[6366 ] = 12'h3a2;
    rom[6367 ] = 12'h3a2;
    rom[6368 ] = 12'h3a2;
    rom[6369 ] = 12'h3a2;
    rom[6370 ] = 12'h3a2;
    rom[6371 ] = 12'h3a2;
    rom[6372 ] = 12'h3a2;
    rom[6373 ] = 12'h3a2;
    rom[6374 ] = 12'h3a2;
    rom[6375 ] = 12'h3a2;
    rom[6376 ] = 12'h3a2;
    rom[6377 ] = 12'h3a2;
    rom[6378 ] = 12'h292;
    rom[6379 ] = 12'h000;
    rom[6380 ] = 12'h000;
    rom[6381 ] = 12'h000;
    rom[6382 ] = 12'h000;
    rom[6383 ] = 12'h000;
    rom[6384 ] = 12'h000;
    rom[6385 ] = 12'h000;
    rom[6386 ] = 12'h000;
    rom[6387 ] = 12'h000;
    rom[6388 ] = 12'h000;
    rom[6389 ] = 12'h000;
    rom[6390 ] = 12'h000;
    rom[6391 ] = 12'h000;
    rom[6392 ] = 12'h000;
    rom[6393 ] = 12'h000;
    rom[6394 ] = 12'h000;
    rom[6395 ] = 12'h000;
    rom[6396 ] = 12'h000;
    rom[6397 ] = 12'h000;
    rom[6398 ] = 12'h000;
    rom[6399 ] = 12'h000;
    rom[6400 ] = 12'h000;
    rom[6401 ] = 12'h5c8;
    rom[6402 ] = 12'h5c8;
    rom[6403 ] = 12'h5c8;
    rom[6404 ] = 12'h5c8;
    rom[6405 ] = 12'h6c7;
    rom[6406 ] = 12'h6c7;
    rom[6407 ] = 12'h6c7;
    rom[6408 ] = 12'h6c7;
    rom[6409 ] = 12'h6c7;
    rom[6410 ] = 12'h6c7;
    rom[6411 ] = 12'h6c7;
    rom[6412 ] = 12'h6c7;
    rom[6413 ] = 12'h6c7;
    rom[6414 ] = 12'h6c7;
    rom[6415 ] = 12'h7c7;
    rom[6416 ] = 12'h7c7;
    rom[6417 ] = 12'h000;
    rom[6418 ] = 12'h000;
    rom[6419 ] = 12'h000;
    rom[6420 ] = 12'h000;
    rom[6421 ] = 12'h000;
    rom[6422 ] = 12'h000;
    rom[6423 ] = 12'h000;
    rom[6424 ] = 12'h000;
    rom[6425 ] = 12'h000;
    rom[6426 ] = 12'h000;
    rom[6427 ] = 12'h000;
    rom[6428 ] = 12'h000;
    rom[6429 ] = 12'h000;
    rom[6430 ] = 12'h000;
    rom[6431 ] = 12'h000;
    rom[6432 ] = 12'h000;
    rom[6433 ] = 12'h000;
    rom[6434 ] = 12'h000;
    rom[6435 ] = 12'h000;
    rom[6436 ] = 12'h000;
    rom[6437 ] = 12'h000;
    rom[6438 ] = 12'h000;
    rom[6439 ] = 12'h492;
    rom[6440 ] = 12'h3a2;
    rom[6441 ] = 12'h3a2;
    rom[6442 ] = 12'h3a2;
    rom[6443 ] = 12'h3a2;
    rom[6444 ] = 12'h3a2;
    rom[6445 ] = 12'h880;
    rom[6446 ] = 12'h000;
    rom[6447 ] = 12'h000;
    rom[6448 ] = 12'h000;
    rom[6449 ] = 12'h000;
    rom[6450 ] = 12'h000;
    rom[6451 ] = 12'h000;
    rom[6452 ] = 12'h000;
    rom[6453 ] = 12'h000;
    rom[6454 ] = 12'h000;
    rom[6455 ] = 12'h000;
    rom[6456 ] = 12'h000;
    rom[6457 ] = 12'h000;
    rom[6458 ] = 12'h000;
    rom[6459 ] = 12'h000;
    rom[6460 ] = 12'h000;
    rom[6461 ] = 12'h000;
    rom[6462 ] = 12'h000;
    rom[6463 ] = 12'h000;
    rom[6464 ] = 12'h000;
    rom[6465 ] = 12'h000;
    rom[6466 ] = 12'h000;
    rom[6467 ] = 12'h000;
    rom[6468 ] = 12'h000;
    rom[6469 ] = 12'h000;
    rom[6470 ] = 12'h000;
    rom[6471 ] = 12'h000;
    rom[6472 ] = 12'h000;
    rom[6473 ] = 12'h000;
    rom[6474 ] = 12'h000;
    rom[6475 ] = 12'h000;
    rom[6476 ] = 12'h000;
    rom[6477 ] = 12'h000;
    rom[6478 ] = 12'h000;
    rom[6479 ] = 12'h000;
    rom[6480 ] = 12'h3a2;
    rom[6481 ] = 12'h3a2;
    rom[6482 ] = 12'h3a2;
    rom[6483 ] = 12'h3a2;
    rom[6484 ] = 12'h3a2;
    rom[6485 ] = 12'h3a2;
    rom[6486 ] = 12'h3a2;
    rom[6487 ] = 12'h3a2;
    rom[6488 ] = 12'h3a2;
    rom[6489 ] = 12'h3a2;
    rom[6490 ] = 12'h3a2;
    rom[6491 ] = 12'h3a2;
    rom[6492 ] = 12'h3a2;
    rom[6493 ] = 12'h3a2;
    rom[6494 ] = 12'h3a2;
    rom[6495 ] = 12'h3a2;
    rom[6496 ] = 12'h3a2;
    rom[6497 ] = 12'h3a2;
    rom[6498 ] = 12'h3a2;
    rom[6499 ] = 12'h3a2;
    rom[6500 ] = 12'h3a2;
    rom[6501 ] = 12'h3a2;
    rom[6502 ] = 12'h3a2;
    rom[6503 ] = 12'h3a2;
    rom[6504 ] = 12'h3a2;
    rom[6505 ] = 12'h000;
    rom[6506 ] = 12'h000;
    rom[6507 ] = 12'h000;
    rom[6508 ] = 12'h000;
    rom[6509 ] = 12'h000;
    rom[6510 ] = 12'h000;
    rom[6511 ] = 12'h000;
    rom[6512 ] = 12'h000;
    rom[6513 ] = 12'h000;
    rom[6514 ] = 12'h000;
    rom[6515 ] = 12'h000;
    rom[6516 ] = 12'h000;
    rom[6517 ] = 12'h000;
    rom[6518 ] = 12'h000;
    rom[6519 ] = 12'h000;
    rom[6520 ] = 12'h000;
    rom[6521 ] = 12'h000;
    rom[6522 ] = 12'h000;
    rom[6523 ] = 12'h000;
    rom[6524 ] = 12'h000;
    rom[6525 ] = 12'h000;
    rom[6526 ] = 12'h000;
    rom[6527 ] = 12'h000;
    rom[6528 ] = 12'h000;
    rom[6529 ] = 12'h5c8;
    rom[6530 ] = 12'h5c8;
    rom[6531 ] = 12'h5c8;
    rom[6532 ] = 12'h5c8;
    rom[6533 ] = 12'h5c8;
    rom[6534 ] = 12'h5c8;
    rom[6535 ] = 12'h6c8;
    rom[6536 ] = 12'h6c7;
    rom[6537 ] = 12'h6c7;
    rom[6538 ] = 12'h6c7;
    rom[6539 ] = 12'h6c7;
    rom[6540 ] = 12'h6c7;
    rom[6541 ] = 12'h6c7;
    rom[6542 ] = 12'h6c7;
    rom[6543 ] = 12'h6c7;
    rom[6544 ] = 12'h696;
    rom[6545 ] = 12'h000;
    rom[6546 ] = 12'h000;
    rom[6547 ] = 12'h000;
    rom[6548 ] = 12'h000;
    rom[6549 ] = 12'h000;
    rom[6550 ] = 12'h000;
    rom[6551 ] = 12'h000;
    rom[6552 ] = 12'h000;
    rom[6553 ] = 12'h000;
    rom[6554 ] = 12'h000;
    rom[6555 ] = 12'h000;
    rom[6556 ] = 12'h000;
    rom[6557 ] = 12'h000;
    rom[6558 ] = 12'h000;
    rom[6559 ] = 12'h000;
    rom[6560 ] = 12'h000;
    rom[6561 ] = 12'h000;
    rom[6562 ] = 12'h000;
    rom[6563 ] = 12'h000;
    rom[6564 ] = 12'h000;
    rom[6565 ] = 12'h000;
    rom[6566 ] = 12'h000;
    rom[6567 ] = 12'h492;
    rom[6568 ] = 12'h3a2;
    rom[6569 ] = 12'h3a2;
    rom[6570 ] = 12'h3a2;
    rom[6571 ] = 12'h3a2;
    rom[6572 ] = 12'h3a2;
    rom[6573 ] = 12'h3a2;
    rom[6574 ] = 12'h3a2;
    rom[6575 ] = 12'h000;
    rom[6576 ] = 12'h000;
    rom[6577 ] = 12'h000;
    rom[6578 ] = 12'h000;
    rom[6579 ] = 12'h000;
    rom[6580 ] = 12'h000;
    rom[6581 ] = 12'h000;
    rom[6582 ] = 12'h000;
    rom[6583 ] = 12'h000;
    rom[6584 ] = 12'h000;
    rom[6585 ] = 12'h000;
    rom[6586 ] = 12'h000;
    rom[6587 ] = 12'h000;
    rom[6588 ] = 12'h000;
    rom[6589 ] = 12'h000;
    rom[6590 ] = 12'h000;
    rom[6591 ] = 12'h000;
    rom[6592 ] = 12'h000;
    rom[6593 ] = 12'h000;
    rom[6594 ] = 12'h000;
    rom[6595 ] = 12'h000;
    rom[6596 ] = 12'h000;
    rom[6597 ] = 12'h000;
    rom[6598 ] = 12'h000;
    rom[6599 ] = 12'h000;
    rom[6600 ] = 12'h000;
    rom[6601 ] = 12'h000;
    rom[6602 ] = 12'h000;
    rom[6603 ] = 12'h000;
    rom[6604 ] = 12'h000;
    rom[6605 ] = 12'h000;
    rom[6606 ] = 12'h3a2;
    rom[6607 ] = 12'h3a2;
    rom[6608 ] = 12'h3a2;
    rom[6609 ] = 12'h3a2;
    rom[6610 ] = 12'h3a2;
    rom[6611 ] = 12'h3a2;
    rom[6612 ] = 12'h3a2;
    rom[6613 ] = 12'h3a2;
    rom[6614 ] = 12'h3a2;
    rom[6615 ] = 12'h3a2;
    rom[6616 ] = 12'h3a2;
    rom[6617 ] = 12'h3a2;
    rom[6618 ] = 12'h3a2;
    rom[6619 ] = 12'h3a2;
    rom[6620 ] = 12'h3a2;
    rom[6621 ] = 12'h3a2;
    rom[6622 ] = 12'h3a2;
    rom[6623 ] = 12'h3a2;
    rom[6624 ] = 12'h3a2;
    rom[6625 ] = 12'h3a2;
    rom[6626 ] = 12'h3a2;
    rom[6627 ] = 12'h3a2;
    rom[6628 ] = 12'h3a2;
    rom[6629 ] = 12'h3a2;
    rom[6630 ] = 12'h3a2;
    rom[6631 ] = 12'h3a2;
    rom[6632 ] = 12'h000;
    rom[6633 ] = 12'h000;
    rom[6634 ] = 12'h000;
    rom[6635 ] = 12'h000;
    rom[6636 ] = 12'h000;
    rom[6637 ] = 12'h000;
    rom[6638 ] = 12'h000;
    rom[6639 ] = 12'h000;
    rom[6640 ] = 12'h000;
    rom[6641 ] = 12'h000;
    rom[6642 ] = 12'h000;
    rom[6643 ] = 12'h000;
    rom[6644 ] = 12'h000;
    rom[6645 ] = 12'h000;
    rom[6646 ] = 12'h000;
    rom[6647 ] = 12'h000;
    rom[6648 ] = 12'h000;
    rom[6649 ] = 12'h000;
    rom[6650 ] = 12'h000;
    rom[6651 ] = 12'h000;
    rom[6652 ] = 12'h000;
    rom[6653 ] = 12'h000;
    rom[6654 ] = 12'h000;
    rom[6655 ] = 12'h000;
    rom[6656 ] = 12'h000;
    rom[6657 ] = 12'h5c8;
    rom[6658 ] = 12'h5c8;
    rom[6659 ] = 12'h5c8;
    rom[6660 ] = 12'h5c8;
    rom[6661 ] = 12'h5c8;
    rom[6662 ] = 12'h5c8;
    rom[6663 ] = 12'h5c8;
    rom[6664 ] = 12'h5c8;
    rom[6665 ] = 12'h5c8;
    rom[6666 ] = 12'h6c7;
    rom[6667 ] = 12'h6c7;
    rom[6668 ] = 12'h6c7;
    rom[6669 ] = 12'h6c7;
    rom[6670 ] = 12'h6c7;
    rom[6671 ] = 12'h6c7;
    rom[6672 ] = 12'h000;
    rom[6673 ] = 12'h000;
    rom[6674 ] = 12'h000;
    rom[6675 ] = 12'h000;
    rom[6676 ] = 12'h000;
    rom[6677 ] = 12'h000;
    rom[6678 ] = 12'h000;
    rom[6679 ] = 12'h000;
    rom[6680 ] = 12'h000;
    rom[6681 ] = 12'h000;
    rom[6682 ] = 12'h000;
    rom[6683 ] = 12'h000;
    rom[6684 ] = 12'h000;
    rom[6685 ] = 12'h000;
    rom[6686 ] = 12'h000;
    rom[6687 ] = 12'h000;
    rom[6688 ] = 12'h000;
    rom[6689 ] = 12'h000;
    rom[6690 ] = 12'h000;
    rom[6691 ] = 12'h000;
    rom[6692 ] = 12'h000;
    rom[6693 ] = 12'h000;
    rom[6694 ] = 12'h000;
    rom[6695 ] = 12'h492;
    rom[6696 ] = 12'h3a2;
    rom[6697 ] = 12'h3a2;
    rom[6698 ] = 12'h3a2;
    rom[6699 ] = 12'h3a2;
    rom[6700 ] = 12'h3a2;
    rom[6701 ] = 12'h3a2;
    rom[6702 ] = 12'h3a2;
    rom[6703 ] = 12'h3a2;
    rom[6704 ] = 12'h3a2;
    rom[6705 ] = 12'h000;
    rom[6706 ] = 12'h000;
    rom[6707 ] = 12'h000;
    rom[6708 ] = 12'h000;
    rom[6709 ] = 12'h000;
    rom[6710 ] = 12'h000;
    rom[6711 ] = 12'h000;
    rom[6712 ] = 12'h000;
    rom[6713 ] = 12'h000;
    rom[6714 ] = 12'h000;
    rom[6715 ] = 12'h000;
    rom[6716 ] = 12'h000;
    rom[6717 ] = 12'h000;
    rom[6718 ] = 12'h000;
    rom[6719 ] = 12'h000;
    rom[6720 ] = 12'h000;
    rom[6721 ] = 12'h000;
    rom[6722 ] = 12'h000;
    rom[6723 ] = 12'h000;
    rom[6724 ] = 12'h000;
    rom[6725 ] = 12'h000;
    rom[6726 ] = 12'h000;
    rom[6727 ] = 12'h000;
    rom[6728 ] = 12'h000;
    rom[6729 ] = 12'h000;
    rom[6730 ] = 12'h000;
    rom[6731 ] = 12'h000;
    rom[6732 ] = 12'h000;
    rom[6733 ] = 12'h3a2;
    rom[6734 ] = 12'h3a2;
    rom[6735 ] = 12'h3a2;
    rom[6736 ] = 12'h3a2;
    rom[6737 ] = 12'h3a2;
    rom[6738 ] = 12'h3a2;
    rom[6739 ] = 12'h3a2;
    rom[6740 ] = 12'h3a2;
    rom[6741 ] = 12'h3a2;
    rom[6742 ] = 12'h3a2;
    rom[6743 ] = 12'h3a2;
    rom[6744 ] = 12'h3a2;
    rom[6745 ] = 12'h3a2;
    rom[6746 ] = 12'h3a2;
    rom[6747 ] = 12'h3a2;
    rom[6748 ] = 12'h3a2;
    rom[6749 ] = 12'h3a2;
    rom[6750 ] = 12'h3a2;
    rom[6751 ] = 12'h3a2;
    rom[6752 ] = 12'h3a2;
    rom[6753 ] = 12'h3a2;
    rom[6754 ] = 12'h3a2;
    rom[6755 ] = 12'h3a2;
    rom[6756 ] = 12'h3a2;
    rom[6757 ] = 12'h3a2;
    rom[6758 ] = 12'h080;
    rom[6759 ] = 12'h000;
    rom[6760 ] = 12'h000;
    rom[6761 ] = 12'h000;
    rom[6762 ] = 12'h000;
    rom[6763 ] = 12'h000;
    rom[6764 ] = 12'h000;
    rom[6765 ] = 12'h000;
    rom[6766 ] = 12'h000;
    rom[6767 ] = 12'h000;
    rom[6768 ] = 12'h000;
    rom[6769 ] = 12'h000;
    rom[6770 ] = 12'h000;
    rom[6771 ] = 12'h000;
    rom[6772 ] = 12'h000;
    rom[6773 ] = 12'h000;
    rom[6774 ] = 12'h000;
    rom[6775 ] = 12'h000;
    rom[6776 ] = 12'h000;
    rom[6777 ] = 12'h000;
    rom[6778 ] = 12'h000;
    rom[6779 ] = 12'h000;
    rom[6780 ] = 12'h000;
    rom[6781 ] = 12'h000;
    rom[6782 ] = 12'h000;
    rom[6783 ] = 12'h000;
    rom[6784 ] = 12'h000;
    rom[6785 ] = 12'h4c9;
    rom[6786 ] = 12'h5c8;
    rom[6787 ] = 12'h5c8;
    rom[6788 ] = 12'h5c8;
    rom[6789 ] = 12'h5c8;
    rom[6790 ] = 12'h5c8;
    rom[6791 ] = 12'h5c8;
    rom[6792 ] = 12'h5c8;
    rom[6793 ] = 12'h5c8;
    rom[6794 ] = 12'h5c8;
    rom[6795 ] = 12'h5c8;
    rom[6796 ] = 12'h6c8;
    rom[6797 ] = 12'h6c7;
    rom[6798 ] = 12'h6c7;
    rom[6799 ] = 12'h6c7;
    rom[6800 ] = 12'h000;
    rom[6801 ] = 12'h000;
    rom[6802 ] = 12'h000;
    rom[6803 ] = 12'h000;
    rom[6804 ] = 12'h000;
    rom[6805 ] = 12'h000;
    rom[6806 ] = 12'h000;
    rom[6807 ] = 12'h000;
    rom[6808 ] = 12'h000;
    rom[6809 ] = 12'h000;
    rom[6810 ] = 12'h000;
    rom[6811 ] = 12'h000;
    rom[6812 ] = 12'h000;
    rom[6813 ] = 12'h000;
    rom[6814 ] = 12'h000;
    rom[6815 ] = 12'h000;
    rom[6816 ] = 12'h000;
    rom[6817 ] = 12'h000;
    rom[6818 ] = 12'h000;
    rom[6819 ] = 12'h000;
    rom[6820 ] = 12'h000;
    rom[6821 ] = 12'h000;
    rom[6822 ] = 12'h000;
    rom[6823 ] = 12'h492;
    rom[6824 ] = 12'h3a2;
    rom[6825 ] = 12'h3a2;
    rom[6826 ] = 12'h3a2;
    rom[6827 ] = 12'h3a2;
    rom[6828 ] = 12'h3a2;
    rom[6829 ] = 12'h3a2;
    rom[6830 ] = 12'h3a2;
    rom[6831 ] = 12'h3a2;
    rom[6832 ] = 12'h3a2;
    rom[6833 ] = 12'h3a2;
    rom[6834 ] = 12'h000;
    rom[6835 ] = 12'h000;
    rom[6836 ] = 12'h000;
    rom[6837 ] = 12'h000;
    rom[6838 ] = 12'h000;
    rom[6839 ] = 12'h000;
    rom[6840 ] = 12'h000;
    rom[6841 ] = 12'h000;
    rom[6842 ] = 12'h000;
    rom[6843 ] = 12'h000;
    rom[6844 ] = 12'h000;
    rom[6845 ] = 12'h000;
    rom[6846 ] = 12'h000;
    rom[6847 ] = 12'h000;
    rom[6848 ] = 12'h000;
    rom[6849 ] = 12'h000;
    rom[6850 ] = 12'h000;
    rom[6851 ] = 12'h000;
    rom[6852 ] = 12'h000;
    rom[6853 ] = 12'h000;
    rom[6854 ] = 12'h000;
    rom[6855 ] = 12'h000;
    rom[6856 ] = 12'h000;
    rom[6857 ] = 12'h000;
    rom[6858 ] = 12'h000;
    rom[6859 ] = 12'h000;
    rom[6860 ] = 12'h3a2;
    rom[6861 ] = 12'h3a2;
    rom[6862 ] = 12'h3a2;
    rom[6863 ] = 12'h3a2;
    rom[6864 ] = 12'h3a2;
    rom[6865 ] = 12'h3a2;
    rom[6866 ] = 12'h3a2;
    rom[6867 ] = 12'h3a2;
    rom[6868 ] = 12'h3a2;
    rom[6869 ] = 12'h3a2;
    rom[6870 ] = 12'h3a2;
    rom[6871 ] = 12'h3a2;
    rom[6872 ] = 12'h3a2;
    rom[6873 ] = 12'h3a2;
    rom[6874 ] = 12'h3a2;
    rom[6875 ] = 12'h3a2;
    rom[6876 ] = 12'h3a2;
    rom[6877 ] = 12'h3a2;
    rom[6878 ] = 12'h3a2;
    rom[6879 ] = 12'h3a2;
    rom[6880 ] = 12'h3a2;
    rom[6881 ] = 12'h3a2;
    rom[6882 ] = 12'h3a2;
    rom[6883 ] = 12'h3a2;
    rom[6884 ] = 12'h3a2;
    rom[6885 ] = 12'h000;
    rom[6886 ] = 12'h000;
    rom[6887 ] = 12'h000;
    rom[6888 ] = 12'h000;
    rom[6889 ] = 12'h000;
    rom[6890 ] = 12'h000;
    rom[6891 ] = 12'h000;
    rom[6892 ] = 12'h000;
    rom[6893 ] = 12'h000;
    rom[6894 ] = 12'h000;
    rom[6895 ] = 12'h000;
    rom[6896 ] = 12'h000;
    rom[6897 ] = 12'h000;
    rom[6898 ] = 12'h000;
    rom[6899 ] = 12'h000;
    rom[6900 ] = 12'h000;
    rom[6901 ] = 12'h000;
    rom[6902 ] = 12'h000;
    rom[6903 ] = 12'h000;
    rom[6904 ] = 12'h000;
    rom[6905 ] = 12'h000;
    rom[6906 ] = 12'h000;
    rom[6907 ] = 12'h000;
    rom[6908 ] = 12'h000;
    rom[6909 ] = 12'h0f0;
    rom[6910 ] = 12'h3a2;
    rom[6911 ] = 12'h000;
    rom[6912 ] = 12'h000;
    rom[6913 ] = 12'h4c9;
    rom[6914 ] = 12'h4c9;
    rom[6915 ] = 12'h4c9;
    rom[6916 ] = 12'h4c8;
    rom[6917 ] = 12'h5c8;
    rom[6918 ] = 12'h5c8;
    rom[6919 ] = 12'h5c8;
    rom[6920 ] = 12'h5c8;
    rom[6921 ] = 12'h5c8;
    rom[6922 ] = 12'h5c8;
    rom[6923 ] = 12'h5c8;
    rom[6924 ] = 12'h5c8;
    rom[6925 ] = 12'h5c8;
    rom[6926 ] = 12'h5c8;
    rom[6927 ] = 12'h6c8;
    rom[6928 ] = 12'h000;
    rom[6929 ] = 12'h000;
    rom[6930 ] = 12'h000;
    rom[6931 ] = 12'h000;
    rom[6932 ] = 12'h000;
    rom[6933 ] = 12'h000;
    rom[6934 ] = 12'h000;
    rom[6935 ] = 12'h000;
    rom[6936 ] = 12'h000;
    rom[6937 ] = 12'h000;
    rom[6938 ] = 12'h000;
    rom[6939 ] = 12'h000;
    rom[6940 ] = 12'h000;
    rom[6941 ] = 12'h000;
    rom[6942 ] = 12'h000;
    rom[6943 ] = 12'h000;
    rom[6944 ] = 12'h000;
    rom[6945 ] = 12'h000;
    rom[6946 ] = 12'h000;
    rom[6947 ] = 12'h000;
    rom[6948 ] = 12'h000;
    rom[6949 ] = 12'h000;
    rom[6950 ] = 12'h000;
    rom[6951 ] = 12'h492;
    rom[6952 ] = 12'h3a2;
    rom[6953 ] = 12'h3a2;
    rom[6954 ] = 12'h3a2;
    rom[6955 ] = 12'h3a2;
    rom[6956 ] = 12'h3a2;
    rom[6957 ] = 12'h3a2;
    rom[6958 ] = 12'h3a2;
    rom[6959 ] = 12'h3a2;
    rom[6960 ] = 12'h3a2;
    rom[6961 ] = 12'h3a2;
    rom[6962 ] = 12'h3a2;
    rom[6963 ] = 12'h3a2;
    rom[6964 ] = 12'h000;
    rom[6965 ] = 12'h000;
    rom[6966 ] = 12'h000;
    rom[6967 ] = 12'h000;
    rom[6968 ] = 12'h000;
    rom[6969 ] = 12'h000;
    rom[6970 ] = 12'h000;
    rom[6971 ] = 12'h000;
    rom[6972 ] = 12'h000;
    rom[6973 ] = 12'h000;
    rom[6974 ] = 12'h000;
    rom[6975 ] = 12'h000;
    rom[6976 ] = 12'h000;
    rom[6977 ] = 12'h000;
    rom[6978 ] = 12'h000;
    rom[6979 ] = 12'h000;
    rom[6980 ] = 12'h000;
    rom[6981 ] = 12'h000;
    rom[6982 ] = 12'h000;
    rom[6983 ] = 12'h000;
    rom[6984 ] = 12'h000;
    rom[6985 ] = 12'h000;
    rom[6986 ] = 12'h3a2;
    rom[6987 ] = 12'h3a2;
    rom[6988 ] = 12'h3a2;
    rom[6989 ] = 12'h3a2;
    rom[6990 ] = 12'h3a2;
    rom[6991 ] = 12'h3a2;
    rom[6992 ] = 12'h3a2;
    rom[6993 ] = 12'h3a2;
    rom[6994 ] = 12'h3a2;
    rom[6995 ] = 12'h3a2;
    rom[6996 ] = 12'h3a2;
    rom[6997 ] = 12'h3a2;
    rom[6998 ] = 12'h3a2;
    rom[6999 ] = 12'h3a2;
    rom[7000 ] = 12'h3a2;
    rom[7001 ] = 12'h3a2;
    rom[7002 ] = 12'h3a2;
    rom[7003 ] = 12'h3a2;
    rom[7004 ] = 12'h3a2;
    rom[7005 ] = 12'h3a2;
    rom[7006 ] = 12'h3a2;
    rom[7007 ] = 12'h3a2;
    rom[7008 ] = 12'h3a2;
    rom[7009 ] = 12'h3a2;
    rom[7010 ] = 12'h3a2;
    rom[7011 ] = 12'h3a2;
    rom[7012 ] = 12'h000;
    rom[7013 ] = 12'h000;
    rom[7014 ] = 12'h000;
    rom[7015 ] = 12'h000;
    rom[7016 ] = 12'h000;
    rom[7017 ] = 12'h000;
    rom[7018 ] = 12'h000;
    rom[7019 ] = 12'h000;
    rom[7020 ] = 12'h000;
    rom[7021 ] = 12'h000;
    rom[7022 ] = 12'h000;
    rom[7023 ] = 12'h000;
    rom[7024 ] = 12'h000;
    rom[7025 ] = 12'h000;
    rom[7026 ] = 12'h000;
    rom[7027 ] = 12'h000;
    rom[7028 ] = 12'h000;
    rom[7029 ] = 12'h000;
    rom[7030 ] = 12'h000;
    rom[7031 ] = 12'h000;
    rom[7032 ] = 12'h000;
    rom[7033 ] = 12'h000;
    rom[7034 ] = 12'h000;
    rom[7035 ] = 12'h000;
    rom[7036 ] = 12'h3a2;
    rom[7037 ] = 12'h3a2;
    rom[7038 ] = 12'h3a2;
    rom[7039 ] = 12'h000;
    rom[7040 ] = 12'h4c9;
    rom[7041 ] = 12'h4c9;
    rom[7042 ] = 12'h4c9;
    rom[7043 ] = 12'h4c9;
    rom[7044 ] = 12'h4c9;
    rom[7045 ] = 12'h4c9;
    rom[7046 ] = 12'h4c9;
    rom[7047 ] = 12'h5c8;
    rom[7048 ] = 12'h5c8;
    rom[7049 ] = 12'h5c8;
    rom[7050 ] = 12'h5c8;
    rom[7051 ] = 12'h5c8;
    rom[7052 ] = 12'h5c8;
    rom[7053 ] = 12'h5c8;
    rom[7054 ] = 12'h5c8;
    rom[7055 ] = 12'h5c8;
    rom[7056 ] = 12'h000;
    rom[7057 ] = 12'h000;
    rom[7058 ] = 12'h000;
    rom[7059 ] = 12'h000;
    rom[7060 ] = 12'h000;
    rom[7061 ] = 12'h000;
    rom[7062 ] = 12'h000;
    rom[7063 ] = 12'h000;
    rom[7064 ] = 12'h000;
    rom[7065 ] = 12'h000;
    rom[7066 ] = 12'h000;
    rom[7067 ] = 12'h000;
    rom[7068 ] = 12'h000;
    rom[7069 ] = 12'h000;
    rom[7070 ] = 12'h000;
    rom[7071 ] = 12'h000;
    rom[7072 ] = 12'h000;
    rom[7073 ] = 12'h000;
    rom[7074 ] = 12'h000;
    rom[7075 ] = 12'h000;
    rom[7076 ] = 12'h000;
    rom[7077 ] = 12'h000;
    rom[7078 ] = 12'h000;
    rom[7079 ] = 12'h492;
    rom[7080 ] = 12'h3a2;
    rom[7081 ] = 12'h3a2;
    rom[7082 ] = 12'h3a2;
    rom[7083 ] = 12'h3a2;
    rom[7084 ] = 12'h3a2;
    rom[7085 ] = 12'h3a2;
    rom[7086 ] = 12'h3a2;
    rom[7087 ] = 12'h3a2;
    rom[7088 ] = 12'h3a2;
    rom[7089 ] = 12'h3a2;
    rom[7090 ] = 12'h3a2;
    rom[7091 ] = 12'h3a2;
    rom[7092 ] = 12'h3a2;
    rom[7093 ] = 12'h000;
    rom[7094 ] = 12'h000;
    rom[7095 ] = 12'h000;
    rom[7096 ] = 12'h000;
    rom[7097 ] = 12'h000;
    rom[7098 ] = 12'h000;
    rom[7099 ] = 12'h000;
    rom[7100 ] = 12'h000;
    rom[7101 ] = 12'h000;
    rom[7102 ] = 12'h000;
    rom[7103 ] = 12'h000;
    rom[7104 ] = 12'h000;
    rom[7105 ] = 12'h000;
    rom[7106 ] = 12'h000;
    rom[7107 ] = 12'h000;
    rom[7108 ] = 12'h000;
    rom[7109 ] = 12'h000;
    rom[7110 ] = 12'h000;
    rom[7111 ] = 12'h000;
    rom[7112 ] = 12'h000;
    rom[7113 ] = 12'h3a2;
    rom[7114 ] = 12'h3a2;
    rom[7115 ] = 12'h3a2;
    rom[7116 ] = 12'h3a2;
    rom[7117 ] = 12'h3a2;
    rom[7118 ] = 12'h3a2;
    rom[7119 ] = 12'h3a2;
    rom[7120 ] = 12'h3a2;
    rom[7121 ] = 12'h3a2;
    rom[7122 ] = 12'h3a2;
    rom[7123 ] = 12'h3a2;
    rom[7124 ] = 12'h3a2;
    rom[7125 ] = 12'h3a2;
    rom[7126 ] = 12'h3a2;
    rom[7127 ] = 12'h3a2;
    rom[7128 ] = 12'h3a2;
    rom[7129 ] = 12'h3a2;
    rom[7130 ] = 12'h3a2;
    rom[7131 ] = 12'h3a2;
    rom[7132 ] = 12'h3a2;
    rom[7133 ] = 12'h3a2;
    rom[7134 ] = 12'h3a2;
    rom[7135 ] = 12'h3a2;
    rom[7136 ] = 12'h3a2;
    rom[7137 ] = 12'h3a2;
    rom[7138 ] = 12'h000;
    rom[7139 ] = 12'h000;
    rom[7140 ] = 12'h000;
    rom[7141 ] = 12'h000;
    rom[7142 ] = 12'h000;
    rom[7143 ] = 12'h000;
    rom[7144 ] = 12'h000;
    rom[7145 ] = 12'h000;
    rom[7146 ] = 12'h000;
    rom[7147 ] = 12'h000;
    rom[7148 ] = 12'h000;
    rom[7149 ] = 12'h000;
    rom[7150 ] = 12'h000;
    rom[7151 ] = 12'h000;
    rom[7152 ] = 12'h000;
    rom[7153 ] = 12'h000;
    rom[7154 ] = 12'h000;
    rom[7155 ] = 12'h000;
    rom[7156 ] = 12'h000;
    rom[7157 ] = 12'h000;
    rom[7158 ] = 12'h000;
    rom[7159 ] = 12'h000;
    rom[7160 ] = 12'h000;
    rom[7161 ] = 12'h000;
    rom[7162 ] = 12'h000;
    rom[7163 ] = 12'h3a2;
    rom[7164 ] = 12'h3a2;
    rom[7165 ] = 12'h3a2;
    rom[7166 ] = 12'h3a2;
    rom[7167 ] = 12'h5a0;
    rom[7168 ] = 12'h4c9;
    rom[7169 ] = 12'h4c9;
    rom[7170 ] = 12'h4c9;
    rom[7171 ] = 12'h4c9;
    rom[7172 ] = 12'h4c9;
    rom[7173 ] = 12'h4c9;
    rom[7174 ] = 12'h4c9;
    rom[7175 ] = 12'h4c9;
    rom[7176 ] = 12'h4c9;
    rom[7177 ] = 12'h4c8;
    rom[7178 ] = 12'h5c8;
    rom[7179 ] = 12'h5c8;
    rom[7180 ] = 12'h5c8;
    rom[7181 ] = 12'h5c8;
    rom[7182 ] = 12'h5c8;
    rom[7183 ] = 12'h000;
    rom[7184 ] = 12'h000;
    rom[7185 ] = 12'h000;
    rom[7186 ] = 12'h000;
    rom[7187 ] = 12'h000;
    rom[7188 ] = 12'h000;
    rom[7189 ] = 12'h000;
    rom[7190 ] = 12'h000;
    rom[7191 ] = 12'h000;
    rom[7192 ] = 12'h000;
    rom[7193 ] = 12'h000;
    rom[7194 ] = 12'h000;
    rom[7195 ] = 12'h000;
    rom[7196 ] = 12'h000;
    rom[7197 ] = 12'h000;
    rom[7198 ] = 12'h000;
    rom[7199 ] = 12'h000;
    rom[7200 ] = 12'h000;
    rom[7201 ] = 12'h000;
    rom[7202 ] = 12'h000;
    rom[7203 ] = 12'h000;
    rom[7204 ] = 12'h000;
    rom[7205 ] = 12'h000;
    rom[7206 ] = 12'h000;
    rom[7207 ] = 12'h492;
    rom[7208 ] = 12'h3a2;
    rom[7209 ] = 12'h3a2;
    rom[7210 ] = 12'h3a2;
    rom[7211 ] = 12'h3a2;
    rom[7212 ] = 12'h3a2;
    rom[7213 ] = 12'h3a2;
    rom[7214 ] = 12'h3a2;
    rom[7215 ] = 12'h3a2;
    rom[7216 ] = 12'h3a2;
    rom[7217 ] = 12'h3a2;
    rom[7218 ] = 12'h3a2;
    rom[7219 ] = 12'h3a2;
    rom[7220 ] = 12'h3a2;
    rom[7221 ] = 12'h3a2;
    rom[7222 ] = 12'h3a2;
    rom[7223 ] = 12'h000;
    rom[7224 ] = 12'h000;
    rom[7225 ] = 12'h000;
    rom[7226 ] = 12'h000;
    rom[7227 ] = 12'h000;
    rom[7228 ] = 12'h000;
    rom[7229 ] = 12'h000;
    rom[7230 ] = 12'h000;
    rom[7231 ] = 12'h000;
    rom[7232 ] = 12'h000;
    rom[7233 ] = 12'h000;
    rom[7234 ] = 12'h000;
    rom[7235 ] = 12'h000;
    rom[7236 ] = 12'h000;
    rom[7237 ] = 12'h000;
    rom[7238 ] = 12'h000;
    rom[7239 ] = 12'h2a1;
    rom[7240 ] = 12'h3a2;
    rom[7241 ] = 12'h3a2;
    rom[7242 ] = 12'h3a2;
    rom[7243 ] = 12'h3a2;
    rom[7244 ] = 12'h3a2;
    rom[7245 ] = 12'h3a2;
    rom[7246 ] = 12'h3a2;
    rom[7247 ] = 12'h3a2;
    rom[7248 ] = 12'h3a2;
    rom[7249 ] = 12'h3a2;
    rom[7250 ] = 12'h3a2;
    rom[7251 ] = 12'h3a2;
    rom[7252 ] = 12'h3a2;
    rom[7253 ] = 12'h3a2;
    rom[7254 ] = 12'h3a2;
    rom[7255 ] = 12'h3a2;
    rom[7256 ] = 12'h3a2;
    rom[7257 ] = 12'h3a2;
    rom[7258 ] = 12'h3a2;
    rom[7259 ] = 12'h3a2;
    rom[7260 ] = 12'h3a2;
    rom[7261 ] = 12'h3a2;
    rom[7262 ] = 12'h3a2;
    rom[7263 ] = 12'h3a2;
    rom[7264 ] = 12'h3a2;
    rom[7265 ] = 12'h000;
    rom[7266 ] = 12'h000;
    rom[7267 ] = 12'h000;
    rom[7268 ] = 12'h000;
    rom[7269 ] = 12'h000;
    rom[7270 ] = 12'h000;
    rom[7271 ] = 12'h000;
    rom[7272 ] = 12'h000;
    rom[7273 ] = 12'h000;
    rom[7274 ] = 12'h000;
    rom[7275 ] = 12'h000;
    rom[7276 ] = 12'h000;
    rom[7277 ] = 12'h000;
    rom[7278 ] = 12'h000;
    rom[7279 ] = 12'h000;
    rom[7280 ] = 12'h000;
    rom[7281 ] = 12'h000;
    rom[7282 ] = 12'h000;
    rom[7283 ] = 12'h000;
    rom[7284 ] = 12'h000;
    rom[7285 ] = 12'h000;
    rom[7286 ] = 12'h000;
    rom[7287 ] = 12'h000;
    rom[7288 ] = 12'h000;
    rom[7289 ] = 12'h0f0;
    rom[7290 ] = 12'h3a2;
    rom[7291 ] = 12'h3a2;
    rom[7292 ] = 12'h3a2;
    rom[7293 ] = 12'h3a2;
    rom[7294 ] = 12'h3a2;
    rom[7295 ] = 12'h3a2;
    rom[7296 ] = 12'h3ca;
    rom[7297 ] = 12'h3c9;
    rom[7298 ] = 12'h4c9;
    rom[7299 ] = 12'h4c9;
    rom[7300 ] = 12'h4c9;
    rom[7301 ] = 12'h4c9;
    rom[7302 ] = 12'h4c9;
    rom[7303 ] = 12'h4c9;
    rom[7304 ] = 12'h4c9;
    rom[7305 ] = 12'h4c9;
    rom[7306 ] = 12'h4c9;
    rom[7307 ] = 12'h4c9;
    rom[7308 ] = 12'h5c8;
    rom[7309 ] = 12'h5c8;
    rom[7310 ] = 12'h5c8;
    rom[7311 ] = 12'h000;
    rom[7312 ] = 12'h000;
    rom[7313 ] = 12'h000;
    rom[7314 ] = 12'h000;
    rom[7315 ] = 12'h000;
    rom[7316 ] = 12'h000;
    rom[7317 ] = 12'h000;
    rom[7318 ] = 12'h000;
    rom[7319 ] = 12'h000;
    rom[7320 ] = 12'h000;
    rom[7321 ] = 12'h000;
    rom[7322 ] = 12'h000;
    rom[7323 ] = 12'h000;
    rom[7324 ] = 12'h000;
    rom[7325 ] = 12'h000;
    rom[7326 ] = 12'h000;
    rom[7327 ] = 12'h000;
    rom[7328 ] = 12'h000;
    rom[7329 ] = 12'h000;
    rom[7330 ] = 12'h000;
    rom[7331 ] = 12'h000;
    rom[7332 ] = 12'h000;
    rom[7333 ] = 12'h000;
    rom[7334 ] = 12'h000;
    rom[7335 ] = 12'h492;
    rom[7336 ] = 12'h3a2;
    rom[7337 ] = 12'h3a2;
    rom[7338 ] = 12'h3a2;
    rom[7339 ] = 12'h3a2;
    rom[7340 ] = 12'h3a2;
    rom[7341 ] = 12'h3a2;
    rom[7342 ] = 12'h3a2;
    rom[7343 ] = 12'h3a2;
    rom[7344 ] = 12'h3a2;
    rom[7345 ] = 12'h3a2;
    rom[7346 ] = 12'h3a2;
    rom[7347 ] = 12'h3a2;
    rom[7348 ] = 12'h3a2;
    rom[7349 ] = 12'h3a2;
    rom[7350 ] = 12'h3a2;
    rom[7351 ] = 12'h3a2;
    rom[7352 ] = 12'h3a2;
    rom[7353 ] = 12'h000;
    rom[7354 ] = 12'h000;
    rom[7355 ] = 12'h000;
    rom[7356 ] = 12'h000;
    rom[7357 ] = 12'h000;
    rom[7358 ] = 12'h000;
    rom[7359 ] = 12'h000;
    rom[7360 ] = 12'h000;
    rom[7361 ] = 12'h000;
    rom[7362 ] = 12'h000;
    rom[7363 ] = 12'h000;
    rom[7364 ] = 12'h000;
    rom[7365 ] = 12'h000;
    rom[7366 ] = 12'h3a2;
    rom[7367 ] = 12'h3a2;
    rom[7368 ] = 12'h3a2;
    rom[7369 ] = 12'h3a2;
    rom[7370 ] = 12'h3a2;
    rom[7371 ] = 12'h3a2;
    rom[7372 ] = 12'h3a2;
    rom[7373 ] = 12'h3a2;
    rom[7374 ] = 12'h3a2;
    rom[7375 ] = 12'h3a2;
    rom[7376 ] = 12'h3a2;
    rom[7377 ] = 12'h3a2;
    rom[7378 ] = 12'h3a2;
    rom[7379 ] = 12'h3a2;
    rom[7380 ] = 12'h3a2;
    rom[7381 ] = 12'h3a2;
    rom[7382 ] = 12'h3a2;
    rom[7383 ] = 12'h3a2;
    rom[7384 ] = 12'h3a2;
    rom[7385 ] = 12'h3a2;
    rom[7386 ] = 12'h3a2;
    rom[7387 ] = 12'h3a2;
    rom[7388 ] = 12'h3a2;
    rom[7389 ] = 12'h3a2;
    rom[7390 ] = 12'h3a2;
    rom[7391 ] = 12'h3a1;
    rom[7392 ] = 12'h000;
    rom[7393 ] = 12'h000;
    rom[7394 ] = 12'h000;
    rom[7395 ] = 12'h000;
    rom[7396 ] = 12'h000;
    rom[7397 ] = 12'h000;
    rom[7398 ] = 12'h000;
    rom[7399 ] = 12'h000;
    rom[7400 ] = 12'h000;
    rom[7401 ] = 12'h000;
    rom[7402 ] = 12'h000;
    rom[7403 ] = 12'h000;
    rom[7404 ] = 12'h000;
    rom[7405 ] = 12'h000;
    rom[7406 ] = 12'h000;
    rom[7407 ] = 12'h000;
    rom[7408 ] = 12'h000;
    rom[7409 ] = 12'h000;
    rom[7410 ] = 12'h000;
    rom[7411 ] = 12'h000;
    rom[7412 ] = 12'h000;
    rom[7413 ] = 12'h000;
    rom[7414 ] = 12'h000;
    rom[7415 ] = 12'h000;
    rom[7416 ] = 12'h3a2;
    rom[7417 ] = 12'h3a2;
    rom[7418 ] = 12'h3a2;
    rom[7419 ] = 12'h3a2;
    rom[7420 ] = 12'h3a2;
    rom[7421 ] = 12'h3a2;
    rom[7422 ] = 12'h3a2;
    rom[7423 ] = 12'h3a2;
    rom[7424 ] = 12'h3ca;
    rom[7425 ] = 12'h3ca;
    rom[7426 ] = 12'h3ca;
    rom[7427 ] = 12'h3c9;
    rom[7428 ] = 12'h3c9;
    rom[7429 ] = 12'h4c9;
    rom[7430 ] = 12'h4c9;
    rom[7431 ] = 12'h4c9;
    rom[7432 ] = 12'h4c9;
    rom[7433 ] = 12'h4c9;
    rom[7434 ] = 12'h4c9;
    rom[7435 ] = 12'h4c9;
    rom[7436 ] = 12'h4c9;
    rom[7437 ] = 12'h4c9;
    rom[7438 ] = 12'h4c9;
    rom[7439 ] = 12'h000;
    rom[7440 ] = 12'h000;
    rom[7441 ] = 12'h000;
    rom[7442 ] = 12'h000;
    rom[7443 ] = 12'h000;
    rom[7444 ] = 12'h000;
    rom[7445 ] = 12'h000;
    rom[7446 ] = 12'h000;
    rom[7447 ] = 12'h000;
    rom[7448 ] = 12'h000;
    rom[7449 ] = 12'h000;
    rom[7450 ] = 12'h000;
    rom[7451 ] = 12'h000;
    rom[7452 ] = 12'h000;
    rom[7453 ] = 12'h000;
    rom[7454 ] = 12'h000;
    rom[7455 ] = 12'h000;
    rom[7456 ] = 12'h000;
    rom[7457 ] = 12'h000;
    rom[7458 ] = 12'h000;
    rom[7459 ] = 12'h000;
    rom[7460 ] = 12'h000;
    rom[7461 ] = 12'h000;
    rom[7462 ] = 12'h000;
    rom[7463 ] = 12'h492;
    rom[7464 ] = 12'h3a2;
    rom[7465 ] = 12'h3a2;
    rom[7466 ] = 12'h3a2;
    rom[7467 ] = 12'h3a2;
    rom[7468 ] = 12'h3a2;
    rom[7469 ] = 12'h3a2;
    rom[7470 ] = 12'h3a2;
    rom[7471 ] = 12'h3a2;
    rom[7472 ] = 12'h3a2;
    rom[7473 ] = 12'h3a2;
    rom[7474 ] = 12'h3a2;
    rom[7475 ] = 12'h3a2;
    rom[7476 ] = 12'h3a2;
    rom[7477 ] = 12'h3a2;
    rom[7478 ] = 12'h3a2;
    rom[7479 ] = 12'h3a2;
    rom[7480 ] = 12'h3a2;
    rom[7481 ] = 12'h3a2;
    rom[7482 ] = 12'h000;
    rom[7483 ] = 12'h000;
    rom[7484 ] = 12'h000;
    rom[7485 ] = 12'h000;
    rom[7486 ] = 12'h000;
    rom[7487 ] = 12'h000;
    rom[7488 ] = 12'h000;
    rom[7489 ] = 12'h000;
    rom[7490 ] = 12'h000;
    rom[7491 ] = 12'h000;
    rom[7492 ] = 12'h000;
    rom[7493 ] = 12'h3a2;
    rom[7494 ] = 12'h3a2;
    rom[7495 ] = 12'h3a2;
    rom[7496 ] = 12'h3a2;
    rom[7497 ] = 12'h3a2;
    rom[7498 ] = 12'h3a2;
    rom[7499 ] = 12'h3a2;
    rom[7500 ] = 12'h3a2;
    rom[7501 ] = 12'h3a2;
    rom[7502 ] = 12'h3a2;
    rom[7503 ] = 12'h3a2;
    rom[7504 ] = 12'h3a2;
    rom[7505 ] = 12'h3a2;
    rom[7506 ] = 12'h3a2;
    rom[7507 ] = 12'h3a2;
    rom[7508 ] = 12'h3a2;
    rom[7509 ] = 12'h3a2;
    rom[7510 ] = 12'h3a2;
    rom[7511 ] = 12'h3a2;
    rom[7512 ] = 12'h3a2;
    rom[7513 ] = 12'h3a2;
    rom[7514 ] = 12'h3a2;
    rom[7515 ] = 12'h3a2;
    rom[7516 ] = 12'h3a2;
    rom[7517 ] = 12'h3a2;
    rom[7518 ] = 12'h000;
    rom[7519 ] = 12'h000;
    rom[7520 ] = 12'h000;
    rom[7521 ] = 12'h000;
    rom[7522 ] = 12'h000;
    rom[7523 ] = 12'h000;
    rom[7524 ] = 12'h000;
    rom[7525 ] = 12'h000;
    rom[7526 ] = 12'h000;
    rom[7527 ] = 12'h000;
    rom[7528 ] = 12'h000;
    rom[7529 ] = 12'h000;
    rom[7530 ] = 12'h000;
    rom[7531 ] = 12'h000;
    rom[7532 ] = 12'h000;
    rom[7533 ] = 12'h000;
    rom[7534 ] = 12'h000;
    rom[7535 ] = 12'h000;
    rom[7536 ] = 12'h000;
    rom[7537 ] = 12'h000;
    rom[7538 ] = 12'h000;
    rom[7539 ] = 12'h000;
    rom[7540 ] = 12'h000;
    rom[7541 ] = 12'h000;
    rom[7542 ] = 12'h000;
    rom[7543 ] = 12'h3a2;
    rom[7544 ] = 12'h3a2;
    rom[7545 ] = 12'h3a2;
    rom[7546 ] = 12'h3a2;
    rom[7547 ] = 12'h3a2;
    rom[7548 ] = 12'h3a2;
    rom[7549 ] = 12'h3a2;
    rom[7550 ] = 12'h3a2;
    rom[7551 ] = 12'h3a2;
    rom[7552 ] = 12'h3ca;
    rom[7553 ] = 12'h3ca;
    rom[7554 ] = 12'h3ca;
    rom[7555 ] = 12'h3ca;
    rom[7556 ] = 12'h3ca;
    rom[7557 ] = 12'h3ca;
    rom[7558 ] = 12'h3c9;
    rom[7559 ] = 12'h4c9;
    rom[7560 ] = 12'h4c9;
    rom[7561 ] = 12'h4c9;
    rom[7562 ] = 12'h4c9;
    rom[7563 ] = 12'h4c9;
    rom[7564 ] = 12'h4c9;
    rom[7565 ] = 12'h4c9;
    rom[7566 ] = 12'h4c9;
    rom[7567 ] = 12'h000;
    rom[7568 ] = 12'h000;
    rom[7569 ] = 12'h000;
    rom[7570 ] = 12'h000;
    rom[7571 ] = 12'h000;
    rom[7572 ] = 12'h000;
    rom[7573 ] = 12'h000;
    rom[7574 ] = 12'h000;
    rom[7575 ] = 12'h000;
    rom[7576 ] = 12'h000;
    rom[7577 ] = 12'h000;
    rom[7578 ] = 12'h000;
    rom[7579 ] = 12'h000;
    rom[7580 ] = 12'h000;
    rom[7581 ] = 12'h000;
    rom[7582 ] = 12'h000;
    rom[7583 ] = 12'h000;
    rom[7584 ] = 12'h000;
    rom[7585 ] = 12'h000;
    rom[7586 ] = 12'h000;
    rom[7587 ] = 12'h000;
    rom[7588 ] = 12'h000;
    rom[7589 ] = 12'h000;
    rom[7590 ] = 12'h000;
    rom[7591 ] = 12'h492;
    rom[7592 ] = 12'h3a2;
    rom[7593 ] = 12'h3a2;
    rom[7594 ] = 12'h3a2;
    rom[7595 ] = 12'h3a2;
    rom[7596 ] = 12'h3a2;
    rom[7597 ] = 12'h3a2;
    rom[7598 ] = 12'h3a2;
    rom[7599 ] = 12'h3a2;
    rom[7600 ] = 12'h3a2;
    rom[7601 ] = 12'h3a2;
    rom[7602 ] = 12'h3a2;
    rom[7603 ] = 12'h3a2;
    rom[7604 ] = 12'h3a2;
    rom[7605 ] = 12'h3a2;
    rom[7606 ] = 12'h3a2;
    rom[7607 ] = 12'h3a2;
    rom[7608 ] = 12'h3a2;
    rom[7609 ] = 12'h3a2;
    rom[7610 ] = 12'h3a2;
    rom[7611 ] = 12'h3a2;
    rom[7612 ] = 12'h000;
    rom[7613 ] = 12'h000;
    rom[7614 ] = 12'h000;
    rom[7615 ] = 12'h000;
    rom[7616 ] = 12'h000;
    rom[7617 ] = 12'h000;
    rom[7618 ] = 12'h000;
    rom[7619 ] = 12'h392;
    rom[7620 ] = 12'h3a2;
    rom[7621 ] = 12'h3a2;
    rom[7622 ] = 12'h3a2;
    rom[7623 ] = 12'h3a2;
    rom[7624 ] = 12'h3a2;
    rom[7625 ] = 12'h3a2;
    rom[7626 ] = 12'h3a2;
    rom[7627 ] = 12'h3a2;
    rom[7628 ] = 12'h3a2;
    rom[7629 ] = 12'h3a2;
    rom[7630 ] = 12'h3a2;
    rom[7631 ] = 12'h3a2;
    rom[7632 ] = 12'h3a2;
    rom[7633 ] = 12'h3a2;
    rom[7634 ] = 12'h3a2;
    rom[7635 ] = 12'h3a2;
    rom[7636 ] = 12'h3a2;
    rom[7637 ] = 12'h3a2;
    rom[7638 ] = 12'h3a2;
    rom[7639 ] = 12'h3a2;
    rom[7640 ] = 12'h3a2;
    rom[7641 ] = 12'h3a2;
    rom[7642 ] = 12'h3a2;
    rom[7643 ] = 12'h3a2;
    rom[7644 ] = 12'h3a2;
    rom[7645 ] = 12'h000;
    rom[7646 ] = 12'h000;
    rom[7647 ] = 12'h000;
    rom[7648 ] = 12'h000;
    rom[7649 ] = 12'h000;
    rom[7650 ] = 12'h000;
    rom[7651 ] = 12'h000;
    rom[7652 ] = 12'h000;
    rom[7653 ] = 12'h000;
    rom[7654 ] = 12'h000;
    rom[7655 ] = 12'h000;
    rom[7656 ] = 12'h000;
    rom[7657 ] = 12'h000;
    rom[7658 ] = 12'h000;
    rom[7659 ] = 12'h000;
    rom[7660 ] = 12'h000;
    rom[7661 ] = 12'h000;
    rom[7662 ] = 12'h000;
    rom[7663 ] = 12'h000;
    rom[7664 ] = 12'h000;
    rom[7665 ] = 12'h000;
    rom[7666 ] = 12'h000;
    rom[7667 ] = 12'h000;
    rom[7668 ] = 12'h000;
    rom[7669 ] = 12'h392;
    rom[7670 ] = 12'h3a2;
    rom[7671 ] = 12'h3a2;
    rom[7672 ] = 12'h3a2;
    rom[7673 ] = 12'h3a2;
    rom[7674 ] = 12'h3a2;
    rom[7675 ] = 12'h3a2;
    rom[7676 ] = 12'h3a2;
    rom[7677 ] = 12'h3a2;
    rom[7678 ] = 12'h3a2;
    rom[7679 ] = 12'h3a2;
    rom[7680 ] = 12'h3ca;
    rom[7681 ] = 12'h3ca;
    rom[7682 ] = 12'h3ca;
    rom[7683 ] = 12'h3ca;
    rom[7684 ] = 12'h3ca;
    rom[7685 ] = 12'h3ca;
    rom[7686 ] = 12'h3ca;
    rom[7687 ] = 12'h3ca;
    rom[7688 ] = 12'h3ca;
    rom[7689 ] = 12'h3c9;
    rom[7690 ] = 12'h4c9;
    rom[7691 ] = 12'h4c9;
    rom[7692 ] = 12'h4c9;
    rom[7693 ] = 12'h4c9;
    rom[7694 ] = 12'h4c9;
    rom[7695 ] = 12'h000;
    rom[7696 ] = 12'h000;
    rom[7697 ] = 12'h000;
    rom[7698 ] = 12'h000;
    rom[7699 ] = 12'h000;
    rom[7700 ] = 12'h000;
    rom[7701 ] = 12'h000;
    rom[7702 ] = 12'h000;
    rom[7703 ] = 12'h000;
    rom[7704 ] = 12'h000;
    rom[7705 ] = 12'h000;
    rom[7706 ] = 12'h000;
    rom[7707 ] = 12'h000;
    rom[7708 ] = 12'h000;
    rom[7709 ] = 12'h000;
    rom[7710 ] = 12'h000;
    rom[7711 ] = 12'h000;
    rom[7712 ] = 12'h000;
    rom[7713 ] = 12'h000;
    rom[7714 ] = 12'h000;
    rom[7715 ] = 12'h000;
    rom[7716 ] = 12'h000;
    rom[7717 ] = 12'h000;
    rom[7718 ] = 12'h000;
    rom[7719 ] = 12'h492;
    rom[7720 ] = 12'h3a2;
    rom[7721 ] = 12'h3a2;
    rom[7722 ] = 12'h3a2;
    rom[7723 ] = 12'h3a2;
    rom[7724 ] = 12'h3a2;
    rom[7725 ] = 12'h3a2;
    rom[7726 ] = 12'h3a2;
    rom[7727 ] = 12'h3a2;
    rom[7728 ] = 12'h3a2;
    rom[7729 ] = 12'h3a2;
    rom[7730 ] = 12'h3a2;
    rom[7731 ] = 12'h3a2;
    rom[7732 ] = 12'h3a2;
    rom[7733 ] = 12'h3a2;
    rom[7734 ] = 12'h3a2;
    rom[7735 ] = 12'h3a2;
    rom[7736 ] = 12'h3a2;
    rom[7737 ] = 12'h3a2;
    rom[7738 ] = 12'h3a2;
    rom[7739 ] = 12'h3a2;
    rom[7740 ] = 12'h3a2;
    rom[7741 ] = 12'h000;
    rom[7742 ] = 12'h000;
    rom[7743 ] = 12'h000;
    rom[7744 ] = 12'h000;
    rom[7745 ] = 12'h000;
    rom[7746 ] = 12'h3a2;
    rom[7747 ] = 12'h3a2;
    rom[7748 ] = 12'h3a2;
    rom[7749 ] = 12'h3a2;
    rom[7750 ] = 12'h3a2;
    rom[7751 ] = 12'h3a2;
    rom[7752 ] = 12'h3a2;
    rom[7753 ] = 12'h3a2;
    rom[7754 ] = 12'h3a2;
    rom[7755 ] = 12'h3a2;
    rom[7756 ] = 12'h3a2;
    rom[7757 ] = 12'h3a2;
    rom[7758 ] = 12'h3a2;
    rom[7759 ] = 12'h3a2;
    rom[7760 ] = 12'h3a2;
    rom[7761 ] = 12'h3a2;
    rom[7762 ] = 12'h3a2;
    rom[7763 ] = 12'h3a2;
    rom[7764 ] = 12'h3a2;
    rom[7765 ] = 12'h3a2;
    rom[7766 ] = 12'h3a2;
    rom[7767 ] = 12'h3a2;
    rom[7768 ] = 12'h3a2;
    rom[7769 ] = 12'h3a2;
    rom[7770 ] = 12'h3a2;
    rom[7771 ] = 12'h392;
    rom[7772 ] = 12'h000;
    rom[7773 ] = 12'h000;
    rom[7774 ] = 12'h000;
    rom[7775 ] = 12'h000;
    rom[7776 ] = 12'h000;
    rom[7777 ] = 12'h000;
    rom[7778 ] = 12'h000;
    rom[7779 ] = 12'h000;
    rom[7780 ] = 12'h000;
    rom[7781 ] = 12'h000;
    rom[7782 ] = 12'h000;
    rom[7783 ] = 12'h000;
    rom[7784 ] = 12'h000;
    rom[7785 ] = 12'h000;
    rom[7786 ] = 12'h000;
    rom[7787 ] = 12'h000;
    rom[7788 ] = 12'h000;
    rom[7789 ] = 12'h000;
    rom[7790 ] = 12'h000;
    rom[7791 ] = 12'h000;
    rom[7792 ] = 12'h000;
    rom[7793 ] = 12'h000;
    rom[7794 ] = 12'h000;
    rom[7795 ] = 12'h000;
    rom[7796 ] = 12'h3a2;
    rom[7797 ] = 12'h3a2;
    rom[7798 ] = 12'h3a2;
    rom[7799 ] = 12'h3a2;
    rom[7800 ] = 12'h3a2;
    rom[7801 ] = 12'h3a2;
    rom[7802 ] = 12'h3a2;
    rom[7803 ] = 12'h3a2;
    rom[7804 ] = 12'h3a2;
    rom[7805 ] = 12'h3a2;
    rom[7806 ] = 12'h3a2;
    rom[7807 ] = 12'h3a2;
    rom[7808 ] = 12'h3ca;
    rom[7809 ] = 12'h3ca;
    rom[7810 ] = 12'h3ca;
    rom[7811 ] = 12'h3ca;
    rom[7812 ] = 12'h3ca;
    rom[7813 ] = 12'h3ca;
    rom[7814 ] = 12'h3ca;
    rom[7815 ] = 12'h3ca;
    rom[7816 ] = 12'h3ca;
    rom[7817 ] = 12'h3ca;
    rom[7818 ] = 12'h3ca;
    rom[7819 ] = 12'h3c9;
    rom[7820 ] = 12'h3c9;
    rom[7821 ] = 12'h4c9;
    rom[7822 ] = 12'h4c9;
    rom[7823 ] = 12'h000;
    rom[7824 ] = 12'h000;
    rom[7825 ] = 12'h000;
    rom[7826 ] = 12'h000;
    rom[7827 ] = 12'h000;
    rom[7828 ] = 12'h000;
    rom[7829 ] = 12'h000;
    rom[7830 ] = 12'h000;
    rom[7831 ] = 12'h000;
    rom[7832 ] = 12'h000;
    rom[7833 ] = 12'h000;
    rom[7834 ] = 12'h000;
    rom[7835 ] = 12'h000;
    rom[7836 ] = 12'h000;
    rom[7837 ] = 12'h000;
    rom[7838 ] = 12'h000;
    rom[7839 ] = 12'h000;
    rom[7840 ] = 12'h000;
    rom[7841 ] = 12'h000;
    rom[7842 ] = 12'h000;
    rom[7843 ] = 12'h000;
    rom[7844 ] = 12'h000;
    rom[7845 ] = 12'h000;
    rom[7846 ] = 12'h000;
    rom[7847 ] = 12'h492;
    rom[7848 ] = 12'h3a2;
    rom[7849 ] = 12'h3a2;
    rom[7850 ] = 12'h3a2;
    rom[7851 ] = 12'h3a2;
    rom[7852 ] = 12'h3a2;
    rom[7853 ] = 12'h3a2;
    rom[7854 ] = 12'h3a2;
    rom[7855 ] = 12'h3a2;
    rom[7856 ] = 12'h3a2;
    rom[7857 ] = 12'h3a2;
    rom[7858 ] = 12'h3a2;
    rom[7859 ] = 12'h3a2;
    rom[7860 ] = 12'h3a2;
    rom[7861 ] = 12'h3a2;
    rom[7862 ] = 12'h3a2;
    rom[7863 ] = 12'h3a2;
    rom[7864 ] = 12'h3a2;
    rom[7865 ] = 12'h3a2;
    rom[7866 ] = 12'h3a2;
    rom[7867 ] = 12'h3a2;
    rom[7868 ] = 12'h3a2;
    rom[7869 ] = 12'h3a2;
    rom[7870 ] = 12'h3a2;
    rom[7871 ] = 12'h000;
    rom[7872 ] = 12'h000;
    rom[7873 ] = 12'h3a2;
    rom[7874 ] = 12'h3a2;
    rom[7875 ] = 12'h3a2;
    rom[7876 ] = 12'h3a2;
    rom[7877 ] = 12'h3a2;
    rom[7878 ] = 12'h3a2;
    rom[7879 ] = 12'h3a2;
    rom[7880 ] = 12'h3a2;
    rom[7881 ] = 12'h3a2;
    rom[7882 ] = 12'h3a2;
    rom[7883 ] = 12'h3a2;
    rom[7884 ] = 12'h3a2;
    rom[7885 ] = 12'h3a2;
    rom[7886 ] = 12'h3a2;
    rom[7887 ] = 12'h3a2;
    rom[7888 ] = 12'h3a2;
    rom[7889 ] = 12'h3a2;
    rom[7890 ] = 12'h3a2;
    rom[7891 ] = 12'h3a2;
    rom[7892 ] = 12'h3a2;
    rom[7893 ] = 12'h3a2;
    rom[7894 ] = 12'h3a2;
    rom[7895 ] = 12'h3a2;
    rom[7896 ] = 12'h3a2;
    rom[7897 ] = 12'h3a2;
    rom[7898 ] = 12'h000;
    rom[7899 ] = 12'h000;
    rom[7900 ] = 12'h000;
    rom[7901 ] = 12'h000;
    rom[7902 ] = 12'h000;
    rom[7903 ] = 12'h000;
    rom[7904 ] = 12'h000;
    rom[7905 ] = 12'h000;
    rom[7906 ] = 12'h000;
    rom[7907 ] = 12'h000;
    rom[7908 ] = 12'h000;
    rom[7909 ] = 12'h000;
    rom[7910 ] = 12'h000;
    rom[7911 ] = 12'h000;
    rom[7912 ] = 12'h000;
    rom[7913 ] = 12'h000;
    rom[7914 ] = 12'h000;
    rom[7915 ] = 12'h000;
    rom[7916 ] = 12'h000;
    rom[7917 ] = 12'h000;
    rom[7918 ] = 12'h000;
    rom[7919 ] = 12'h000;
    rom[7920 ] = 12'h000;
    rom[7921 ] = 12'h000;
    rom[7922 ] = 12'h000;
    rom[7923 ] = 12'h3a2;
    rom[7924 ] = 12'h3a2;
    rom[7925 ] = 12'h3a2;
    rom[7926 ] = 12'h3a2;
    rom[7927 ] = 12'h3a2;
    rom[7928 ] = 12'h3a2;
    rom[7929 ] = 12'h3a2;
    rom[7930 ] = 12'h3a2;
    rom[7931 ] = 12'h3a2;
    rom[7932 ] = 12'h3a2;
    rom[7933 ] = 12'h3a2;
    rom[7934 ] = 12'h3a2;
    rom[7935 ] = 12'h3a2;
    rom[7936 ] = 12'h3ca;
    rom[7937 ] = 12'h3ca;
    rom[7938 ] = 12'h3ca;
    rom[7939 ] = 12'h3ca;
    rom[7940 ] = 12'h3ca;
    rom[7941 ] = 12'h3ca;
    rom[7942 ] = 12'h3ca;
    rom[7943 ] = 12'h3ca;
    rom[7944 ] = 12'h3ca;
    rom[7945 ] = 12'h3ca;
    rom[7946 ] = 12'h3ca;
    rom[7947 ] = 12'h3ca;
    rom[7948 ] = 12'h3ca;
    rom[7949 ] = 12'h3ca;
    rom[7950 ] = 12'h3c9;
    rom[7951 ] = 12'h000;
    rom[7952 ] = 12'h000;
    rom[7953 ] = 12'h000;
    rom[7954 ] = 12'h000;
    rom[7955 ] = 12'h000;
    rom[7956 ] = 12'h000;
    rom[7957 ] = 12'h000;
    rom[7958 ] = 12'h000;
    rom[7959 ] = 12'h000;
    rom[7960 ] = 12'h000;
    rom[7961 ] = 12'h000;
    rom[7962 ] = 12'h000;
    rom[7963 ] = 12'h000;
    rom[7964 ] = 12'h000;
    rom[7965 ] = 12'h000;
    rom[7966 ] = 12'h000;
    rom[7967 ] = 12'h000;
    rom[7968 ] = 12'h000;
    rom[7969 ] = 12'h000;
    rom[7970 ] = 12'h000;
    rom[7971 ] = 12'h000;
    rom[7972 ] = 12'h000;
    rom[7973 ] = 12'h000;
    rom[7974 ] = 12'h000;
    rom[7975 ] = 12'h492;
    rom[7976 ] = 12'h3a2;
    rom[7977 ] = 12'h3a2;
    rom[7978 ] = 12'h3a2;
    rom[7979 ] = 12'h3a2;
    rom[7980 ] = 12'h3a2;
    rom[7981 ] = 12'h3a2;
    rom[7982 ] = 12'h3a2;
    rom[7983 ] = 12'h3a2;
    rom[7984 ] = 12'h3a2;
    rom[7985 ] = 12'h3a2;
    rom[7986 ] = 12'h3a2;
    rom[7987 ] = 12'h3a2;
    rom[7988 ] = 12'h3a2;
    rom[7989 ] = 12'h3a2;
    rom[7990 ] = 12'h3a2;
    rom[7991 ] = 12'h3a2;
    rom[7992 ] = 12'h3a2;
    rom[7993 ] = 12'h3a2;
    rom[7994 ] = 12'h3a2;
    rom[7995 ] = 12'h3a2;
    rom[7996 ] = 12'h3a2;
    rom[7997 ] = 12'h3a2;
    rom[7998 ] = 12'h3a2;
    rom[7999 ] = 12'h3a2;
    rom[8000 ] = 12'h3a2;
    rom[8001 ] = 12'h3a2;
    rom[8002 ] = 12'h3a2;
    rom[8003 ] = 12'h3a2;
    rom[8004 ] = 12'h3a2;
    rom[8005 ] = 12'h3a2;
    rom[8006 ] = 12'h3a2;
    rom[8007 ] = 12'h3a2;
    rom[8008 ] = 12'h3a2;
    rom[8009 ] = 12'h3a2;
    rom[8010 ] = 12'h3a2;
    rom[8011 ] = 12'h3a2;
    rom[8012 ] = 12'h3a2;
    rom[8013 ] = 12'h3a2;
    rom[8014 ] = 12'h3a2;
    rom[8015 ] = 12'h3a2;
    rom[8016 ] = 12'h3a2;
    rom[8017 ] = 12'h3a2;
    rom[8018 ] = 12'h3a2;
    rom[8019 ] = 12'h3a2;
    rom[8020 ] = 12'h3a2;
    rom[8021 ] = 12'h3a2;
    rom[8022 ] = 12'h3a2;
    rom[8023 ] = 12'h3a2;
    rom[8024 ] = 12'h3a2;
    rom[8025 ] = 12'h000;
    rom[8026 ] = 12'h000;
    rom[8027 ] = 12'h000;
    rom[8028 ] = 12'h000;
    rom[8029 ] = 12'h000;
    rom[8030 ] = 12'h000;
    rom[8031 ] = 12'h000;
    rom[8032 ] = 12'h000;
    rom[8033 ] = 12'h000;
    rom[8034 ] = 12'h000;
    rom[8035 ] = 12'h000;
    rom[8036 ] = 12'h000;
    rom[8037 ] = 12'h000;
    rom[8038 ] = 12'h000;
    rom[8039 ] = 12'h000;
    rom[8040 ] = 12'h000;
    rom[8041 ] = 12'h000;
    rom[8042 ] = 12'h000;
    rom[8043 ] = 12'h000;
    rom[8044 ] = 12'h000;
    rom[8045 ] = 12'h000;
    rom[8046 ] = 12'h000;
    rom[8047 ] = 12'h000;
    rom[8048 ] = 12'h000;
    rom[8049 ] = 12'h392;
    rom[8050 ] = 12'h3a2;
    rom[8051 ] = 12'h3a2;
    rom[8052 ] = 12'h3a2;
    rom[8053 ] = 12'h3a2;
    rom[8054 ] = 12'h3a2;
    rom[8055 ] = 12'h3a2;
    rom[8056 ] = 12'h3a2;
    rom[8057 ] = 12'h3a2;
    rom[8058 ] = 12'h3a2;
    rom[8059 ] = 12'h3a2;
    rom[8060 ] = 12'h3a2;
    rom[8061 ] = 12'h3a2;
    rom[8062 ] = 12'h3a2;
    rom[8063 ] = 12'h3a2;
    rom[8064 ] = 12'h3ca;
    rom[8065 ] = 12'h3ca;
    rom[8066 ] = 12'h3ca;
    rom[8067 ] = 12'h3ca;
    rom[8068 ] = 12'h3ca;
    rom[8069 ] = 12'h3ca;
    rom[8070 ] = 12'h3ca;
    rom[8071 ] = 12'h3ca;
    rom[8072 ] = 12'h3ca;
    rom[8073 ] = 12'h3ca;
    rom[8074 ] = 12'h3ca;
    rom[8075 ] = 12'h3ca;
    rom[8076 ] = 12'h3ca;
    rom[8077 ] = 12'h3ca;
    rom[8078 ] = 12'h3ca;
    rom[8079 ] = 12'h000;
    rom[8080 ] = 12'h000;
    rom[8081 ] = 12'h000;
    rom[8082 ] = 12'h000;
    rom[8083 ] = 12'h000;
    rom[8084 ] = 12'h000;
    rom[8085 ] = 12'h000;
    rom[8086 ] = 12'h000;
    rom[8087 ] = 12'h000;
    rom[8088 ] = 12'h000;
    rom[8089 ] = 12'h000;
    rom[8090 ] = 12'h000;
    rom[8091 ] = 12'h000;
    rom[8092 ] = 12'h000;
    rom[8093 ] = 12'h000;
    rom[8094 ] = 12'h000;
    rom[8095 ] = 12'h000;
    rom[8096 ] = 12'h000;
    rom[8097 ] = 12'h000;
    rom[8098 ] = 12'h000;
    rom[8099 ] = 12'h000;
    rom[8100 ] = 12'h000;
    rom[8101 ] = 12'h000;
    rom[8102 ] = 12'h000;
    rom[8103 ] = 12'h492;
    rom[8104 ] = 12'h3a2;
    rom[8105 ] = 12'h3a2;
    rom[8106 ] = 12'h3a2;
    rom[8107 ] = 12'h3a2;
    rom[8108 ] = 12'h3a2;
    rom[8109 ] = 12'h3a2;
    rom[8110 ] = 12'h3a2;
    rom[8111 ] = 12'h3a2;
    rom[8112 ] = 12'h3a2;
    rom[8113 ] = 12'h3a2;
    rom[8114 ] = 12'h3a2;
    rom[8115 ] = 12'h3a2;
    rom[8116 ] = 12'h3a2;
    rom[8117 ] = 12'h3a2;
    rom[8118 ] = 12'h3a2;
    rom[8119 ] = 12'h3a2;
    rom[8120 ] = 12'h3a2;
    rom[8121 ] = 12'h3a2;
    rom[8122 ] = 12'h3a2;
    rom[8123 ] = 12'h3a2;
    rom[8124 ] = 12'h3a2;
    rom[8125 ] = 12'h3a2;
    rom[8126 ] = 12'h3a2;
    rom[8127 ] = 12'h3a2;
    rom[8128 ] = 12'h3a2;
    rom[8129 ] = 12'h3a2;
    rom[8130 ] = 12'h3a2;
    rom[8131 ] = 12'h3a2;
    rom[8132 ] = 12'h3a2;
    rom[8133 ] = 12'h3a2;
    rom[8134 ] = 12'h3a2;
    rom[8135 ] = 12'h3a2;
    rom[8136 ] = 12'h3a2;
    rom[8137 ] = 12'h3a2;
    rom[8138 ] = 12'h3a2;
    rom[8139 ] = 12'h3a2;
    rom[8140 ] = 12'h3a2;
    rom[8141 ] = 12'h3a2;
    rom[8142 ] = 12'h3a2;
    rom[8143 ] = 12'h3a2;
    rom[8144 ] = 12'h3a2;
    rom[8145 ] = 12'h3a2;
    rom[8146 ] = 12'h3a2;
    rom[8147 ] = 12'h3a2;
    rom[8148 ] = 12'h3a2;
    rom[8149 ] = 12'h3a2;
    rom[8150 ] = 12'h3a2;
    rom[8151 ] = 12'h3a1;
    rom[8152 ] = 12'h000;
    rom[8153 ] = 12'h000;
    rom[8154 ] = 12'h000;
    rom[8155 ] = 12'h000;
    rom[8156 ] = 12'h000;
    rom[8157 ] = 12'h000;
    rom[8158 ] = 12'h000;
    rom[8159 ] = 12'h000;
    rom[8160 ] = 12'h000;
    rom[8161 ] = 12'h000;
    rom[8162 ] = 12'h000;
    rom[8163 ] = 12'h000;
    rom[8164 ] = 12'h000;
    rom[8165 ] = 12'h000;
    rom[8166 ] = 12'h000;
    rom[8167 ] = 12'h000;
    rom[8168 ] = 12'h000;
    rom[8169 ] = 12'h000;
    rom[8170 ] = 12'h000;
    rom[8171 ] = 12'h000;
    rom[8172 ] = 12'h000;
    rom[8173 ] = 12'h000;
    rom[8174 ] = 12'h000;
    rom[8175 ] = 12'h000;
    rom[8176 ] = 12'h000;
    rom[8177 ] = 12'h3a2;
    rom[8178 ] = 12'h3a2;
    rom[8179 ] = 12'h3a2;
    rom[8180 ] = 12'h3a2;
    rom[8181 ] = 12'h3a2;
    rom[8182 ] = 12'h3a2;
    rom[8183 ] = 12'h3a2;
    rom[8184 ] = 12'h3a2;
    rom[8185 ] = 12'h3a2;
    rom[8186 ] = 12'h3a2;
    rom[8187 ] = 12'h3a2;
    rom[8188 ] = 12'h3a2;
    rom[8189 ] = 12'h3a2;
    rom[8190 ] = 12'h3a2;
    rom[8191 ] = 12'h3a2;
    rom[8192 ] = 12'h3ca;
    rom[8193 ] = 12'h3ca;
    rom[8194 ] = 12'h3ca;
    rom[8195 ] = 12'h3ca;
    rom[8196 ] = 12'h3ca;
    rom[8197 ] = 12'h3ca;
    rom[8198 ] = 12'h3ca;
    rom[8199 ] = 12'h3ca;
    rom[8200 ] = 12'h3ca;
    rom[8201 ] = 12'h3ca;
    rom[8202 ] = 12'h3ca;
    rom[8203 ] = 12'h3ca;
    rom[8204 ] = 12'h3ca;
    rom[8205 ] = 12'h3ca;
    rom[8206 ] = 12'h3ca;
    rom[8207 ] = 12'h000;
    rom[8208 ] = 12'h000;
    rom[8209 ] = 12'h000;
    rom[8210 ] = 12'h000;
    rom[8211 ] = 12'h000;
    rom[8212 ] = 12'h000;
    rom[8213 ] = 12'h000;
    rom[8214 ] = 12'h000;
    rom[8215 ] = 12'h000;
    rom[8216 ] = 12'h000;
    rom[8217 ] = 12'h000;
    rom[8218 ] = 12'h000;
    rom[8219 ] = 12'h000;
    rom[8220 ] = 12'h000;
    rom[8221 ] = 12'h000;
    rom[8222 ] = 12'h000;
    rom[8223 ] = 12'h000;
    rom[8224 ] = 12'h000;
    rom[8225 ] = 12'h000;
    rom[8226 ] = 12'h000;
    rom[8227 ] = 12'h000;
    rom[8228 ] = 12'h000;
    rom[8229 ] = 12'h000;
    rom[8230 ] = 12'h000;
    rom[8231 ] = 12'h492;
    rom[8232 ] = 12'h3a2;
    rom[8233 ] = 12'h3a2;
    rom[8234 ] = 12'h3a2;
    rom[8235 ] = 12'h3a2;
    rom[8236 ] = 12'h3a2;
    rom[8237 ] = 12'h3a2;
    rom[8238 ] = 12'h3a2;
    rom[8239 ] = 12'h3a2;
    rom[8240 ] = 12'h3a2;
    rom[8241 ] = 12'h3a2;
    rom[8242 ] = 12'h3a2;
    rom[8243 ] = 12'h3a2;
    rom[8244 ] = 12'h3a2;
    rom[8245 ] = 12'h3a2;
    rom[8246 ] = 12'h3a2;
    rom[8247 ] = 12'h3a2;
    rom[8248 ] = 12'h3a2;
    rom[8249 ] = 12'h3a2;
    rom[8250 ] = 12'h3a2;
    rom[8251 ] = 12'h3a2;
    rom[8252 ] = 12'h3a2;
    rom[8253 ] = 12'h3a2;
    rom[8254 ] = 12'h3a2;
    rom[8255 ] = 12'h3a2;
    rom[8256 ] = 12'h3a2;
    rom[8257 ] = 12'h3a2;
    rom[8258 ] = 12'h3a2;
    rom[8259 ] = 12'h3a2;
    rom[8260 ] = 12'h3a2;
    rom[8261 ] = 12'h3a2;
    rom[8262 ] = 12'h3a2;
    rom[8263 ] = 12'h3a2;
    rom[8264 ] = 12'h3a2;
    rom[8265 ] = 12'h3a2;
    rom[8266 ] = 12'h3a2;
    rom[8267 ] = 12'h3a2;
    rom[8268 ] = 12'h3a2;
    rom[8269 ] = 12'h3a2;
    rom[8270 ] = 12'h3a2;
    rom[8271 ] = 12'h3a2;
    rom[8272 ] = 12'h3a2;
    rom[8273 ] = 12'h3a2;
    rom[8274 ] = 12'h3a2;
    rom[8275 ] = 12'h3a2;
    rom[8276 ] = 12'h3a2;
    rom[8277 ] = 12'h3a2;
    rom[8278 ] = 12'h000;
    rom[8279 ] = 12'h000;
    rom[8280 ] = 12'h000;
    rom[8281 ] = 12'h000;
    rom[8282 ] = 12'h000;
    rom[8283 ] = 12'h000;
    rom[8284 ] = 12'h000;
    rom[8285 ] = 12'h000;
    rom[8286 ] = 12'h000;
    rom[8287 ] = 12'h000;
    rom[8288 ] = 12'h000;
    rom[8289 ] = 12'h000;
    rom[8290 ] = 12'h000;
    rom[8291 ] = 12'h000;
    rom[8292 ] = 12'h000;
    rom[8293 ] = 12'h000;
    rom[8294 ] = 12'h000;
    rom[8295 ] = 12'h000;
    rom[8296 ] = 12'h000;
    rom[8297 ] = 12'h000;
    rom[8298 ] = 12'h000;
    rom[8299 ] = 12'h000;
    rom[8300 ] = 12'h000;
    rom[8301 ] = 12'h000;
    rom[8302 ] = 12'h000;
    rom[8303 ] = 12'h000;
    rom[8304 ] = 12'h000;
    rom[8305 ] = 12'h3a2;
    rom[8306 ] = 12'h3a2;
    rom[8307 ] = 12'h3a2;
    rom[8308 ] = 12'h3a2;
    rom[8309 ] = 12'h3a2;
    rom[8310 ] = 12'h3a2;
    rom[8311 ] = 12'h3a2;
    rom[8312 ] = 12'h3a2;
    rom[8313 ] = 12'h3a2;
    rom[8314 ] = 12'h3a2;
    rom[8315 ] = 12'h3a2;
    rom[8316 ] = 12'h3a2;
    rom[8317 ] = 12'h3a2;
    rom[8318 ] = 12'h3a2;
    rom[8319 ] = 12'h3a2;
    rom[8320 ] = 12'h3ca;
    rom[8321 ] = 12'h3ca;
    rom[8322 ] = 12'h3ca;
    rom[8323 ] = 12'h3ca;
    rom[8324 ] = 12'h3ca;
    rom[8325 ] = 12'h3ca;
    rom[8326 ] = 12'h3ca;
    rom[8327 ] = 12'h3ca;
    rom[8328 ] = 12'h3ca;
    rom[8329 ] = 12'h3ca;
    rom[8330 ] = 12'h3ca;
    rom[8331 ] = 12'h3ca;
    rom[8332 ] = 12'h3ca;
    rom[8333 ] = 12'h3ca;
    rom[8334 ] = 12'h3ca;
    rom[8335 ] = 12'h000;
    rom[8336 ] = 12'h000;
    rom[8337 ] = 12'h000;
    rom[8338 ] = 12'h000;
    rom[8339 ] = 12'h000;
    rom[8340 ] = 12'h000;
    rom[8341 ] = 12'h000;
    rom[8342 ] = 12'h000;
    rom[8343 ] = 12'h000;
    rom[8344 ] = 12'h000;
    rom[8345 ] = 12'h000;
    rom[8346 ] = 12'h000;
    rom[8347 ] = 12'h000;
    rom[8348 ] = 12'h000;
    rom[8349 ] = 12'h000;
    rom[8350 ] = 12'h000;
    rom[8351 ] = 12'h000;
    rom[8352 ] = 12'h000;
    rom[8353 ] = 12'h000;
    rom[8354 ] = 12'h000;
    rom[8355 ] = 12'h000;
    rom[8356 ] = 12'h000;
    rom[8357 ] = 12'h000;
    rom[8358 ] = 12'h000;
    rom[8359 ] = 12'h000;
    rom[8360 ] = 12'h3a2;
    rom[8361 ] = 12'h3a2;
    rom[8362 ] = 12'h3a2;
    rom[8363 ] = 12'h3a2;
    rom[8364 ] = 12'h3a2;
    rom[8365 ] = 12'h3a2;
    rom[8366 ] = 12'h3a2;
    rom[8367 ] = 12'h3a2;
    rom[8368 ] = 12'h3a2;
    rom[8369 ] = 12'h3a2;
    rom[8370 ] = 12'h3a2;
    rom[8371 ] = 12'h3a2;
    rom[8372 ] = 12'h3a2;
    rom[8373 ] = 12'h3a2;
    rom[8374 ] = 12'h3a2;
    rom[8375 ] = 12'h3a2;
    rom[8376 ] = 12'h3a2;
    rom[8377 ] = 12'h3a2;
    rom[8378 ] = 12'h3a2;
    rom[8379 ] = 12'h3a2;
    rom[8380 ] = 12'h3a2;
    rom[8381 ] = 12'h3a2;
    rom[8382 ] = 12'h3a2;
    rom[8383 ] = 12'h3a2;
    rom[8384 ] = 12'h3a2;
    rom[8385 ] = 12'h3a2;
    rom[8386 ] = 12'h3a2;
    rom[8387 ] = 12'h3a2;
    rom[8388 ] = 12'h3a2;
    rom[8389 ] = 12'h3a2;
    rom[8390 ] = 12'h3a2;
    rom[8391 ] = 12'h3a2;
    rom[8392 ] = 12'h3a2;
    rom[8393 ] = 12'h3a2;
    rom[8394 ] = 12'h3a2;
    rom[8395 ] = 12'h3a2;
    rom[8396 ] = 12'h3a2;
    rom[8397 ] = 12'h3a2;
    rom[8398 ] = 12'h3a2;
    rom[8399 ] = 12'h3a2;
    rom[8400 ] = 12'h3a2;
    rom[8401 ] = 12'h3a2;
    rom[8402 ] = 12'h3a2;
    rom[8403 ] = 12'h3a2;
    rom[8404 ] = 12'h3a2;
    rom[8405 ] = 12'h000;
    rom[8406 ] = 12'h000;
    rom[8407 ] = 12'h000;
    rom[8408 ] = 12'h000;
    rom[8409 ] = 12'h000;
    rom[8410 ] = 12'h000;
    rom[8411 ] = 12'h000;
    rom[8412 ] = 12'h000;
    rom[8413 ] = 12'h000;
    rom[8414 ] = 12'h000;
    rom[8415 ] = 12'h000;
    rom[8416 ] = 12'h000;
    rom[8417 ] = 12'h000;
    rom[8418 ] = 12'h000;
    rom[8419 ] = 12'h000;
    rom[8420 ] = 12'h000;
    rom[8421 ] = 12'h000;
    rom[8422 ] = 12'h000;
    rom[8423 ] = 12'h000;
    rom[8424 ] = 12'h000;
    rom[8425 ] = 12'h000;
    rom[8426 ] = 12'h000;
    rom[8427 ] = 12'h000;
    rom[8428 ] = 12'h000;
    rom[8429 ] = 12'h000;
    rom[8430 ] = 12'h000;
    rom[8431 ] = 12'h000;
    rom[8432 ] = 12'h000;
    rom[8433 ] = 12'h3a2;
    rom[8434 ] = 12'h3a2;
    rom[8435 ] = 12'h3a2;
    rom[8436 ] = 12'h3a2;
    rom[8437 ] = 12'h3a2;
    rom[8438 ] = 12'h3a2;
    rom[8439 ] = 12'h3a2;
    rom[8440 ] = 12'h3a2;
    rom[8441 ] = 12'h3a2;
    rom[8442 ] = 12'h3a2;
    rom[8443 ] = 12'h3a2;
    rom[8444 ] = 12'h3a2;
    rom[8445 ] = 12'h3a2;
    rom[8446 ] = 12'h3a2;
    rom[8447 ] = 12'h3a2;
    rom[8448 ] = 12'h3ca;
    rom[8449 ] = 12'h3ca;
    rom[8450 ] = 12'h3ca;
    rom[8451 ] = 12'h3ca;
    rom[8452 ] = 12'h3ca;
    rom[8453 ] = 12'h3ca;
    rom[8454 ] = 12'h3ca;
    rom[8455 ] = 12'h3ca;
    rom[8456 ] = 12'h3ca;
    rom[8457 ] = 12'h3ca;
    rom[8458 ] = 12'h3ca;
    rom[8459 ] = 12'h3ca;
    rom[8460 ] = 12'h3ca;
    rom[8461 ] = 12'h3ca;
    rom[8462 ] = 12'h3ca;
    rom[8463 ] = 12'h000;
    rom[8464 ] = 12'h000;
    rom[8465 ] = 12'h000;
    rom[8466 ] = 12'h000;
    rom[8467 ] = 12'h000;
    rom[8468 ] = 12'h000;
    rom[8469 ] = 12'h000;
    rom[8470 ] = 12'h000;
    rom[8471 ] = 12'h000;
    rom[8472 ] = 12'h000;
    rom[8473 ] = 12'h000;
    rom[8474 ] = 12'h000;
    rom[8475 ] = 12'h000;
    rom[8476 ] = 12'h000;
    rom[8477 ] = 12'h000;
    rom[8478 ] = 12'h000;
    rom[8479 ] = 12'h000;
    rom[8480 ] = 12'h000;
    rom[8481 ] = 12'h000;
    rom[8482 ] = 12'h000;
    rom[8483 ] = 12'h000;
    rom[8484 ] = 12'h000;
    rom[8485 ] = 12'h000;
    rom[8486 ] = 12'h000;
    rom[8487 ] = 12'h000;
    rom[8488 ] = 12'h000;
    rom[8489 ] = 12'h392;
    rom[8490 ] = 12'h3a2;
    rom[8491 ] = 12'h3a2;
    rom[8492 ] = 12'h3a2;
    rom[8493 ] = 12'h3a2;
    rom[8494 ] = 12'h3a2;
    rom[8495 ] = 12'h3a2;
    rom[8496 ] = 12'h3a2;
    rom[8497 ] = 12'h3a2;
    rom[8498 ] = 12'h3a2;
    rom[8499 ] = 12'h3a2;
    rom[8500 ] = 12'h3a2;
    rom[8501 ] = 12'h3a2;
    rom[8502 ] = 12'h3a2;
    rom[8503 ] = 12'h3a2;
    rom[8504 ] = 12'h3a2;
    rom[8505 ] = 12'h3a2;
    rom[8506 ] = 12'h3a2;
    rom[8507 ] = 12'h3a2;
    rom[8508 ] = 12'h3a2;
    rom[8509 ] = 12'h3a2;
    rom[8510 ] = 12'h3a2;
    rom[8511 ] = 12'h3a2;
    rom[8512 ] = 12'h3a2;
    rom[8513 ] = 12'h3a2;
    rom[8514 ] = 12'h3a2;
    rom[8515 ] = 12'h3a2;
    rom[8516 ] = 12'h3a2;
    rom[8517 ] = 12'h3a2;
    rom[8518 ] = 12'h3a2;
    rom[8519 ] = 12'h3a2;
    rom[8520 ] = 12'h3a2;
    rom[8521 ] = 12'h3a2;
    rom[8522 ] = 12'h3a2;
    rom[8523 ] = 12'h3a2;
    rom[8524 ] = 12'h3a2;
    rom[8525 ] = 12'h3a2;
    rom[8526 ] = 12'h3a2;
    rom[8527 ] = 12'h3a2;
    rom[8528 ] = 12'h3a2;
    rom[8529 ] = 12'h3a2;
    rom[8530 ] = 12'h3a2;
    rom[8531 ] = 12'h393;
    rom[8532 ] = 12'h000;
    rom[8533 ] = 12'h000;
    rom[8534 ] = 12'h000;
    rom[8535 ] = 12'h000;
    rom[8536 ] = 12'h000;
    rom[8537 ] = 12'h000;
    rom[8538 ] = 12'h000;
    rom[8539 ] = 12'h000;
    rom[8540 ] = 12'h000;
    rom[8541 ] = 12'h000;
    rom[8542 ] = 12'h000;
    rom[8543 ] = 12'h000;
    rom[8544 ] = 12'h000;
    rom[8545 ] = 12'h000;
    rom[8546 ] = 12'h000;
    rom[8547 ] = 12'h000;
    rom[8548 ] = 12'h000;
    rom[8549 ] = 12'h000;
    rom[8550 ] = 12'h000;
    rom[8551 ] = 12'h000;
    rom[8552 ] = 12'h000;
    rom[8553 ] = 12'h000;
    rom[8554 ] = 12'h000;
    rom[8555 ] = 12'h000;
    rom[8556 ] = 12'h000;
    rom[8557 ] = 12'h000;
    rom[8558 ] = 12'h000;
    rom[8559 ] = 12'h000;
    rom[8560 ] = 12'h000;
    rom[8561 ] = 12'h3a2;
    rom[8562 ] = 12'h3a2;
    rom[8563 ] = 12'h3a2;
    rom[8564 ] = 12'h3a2;
    rom[8565 ] = 12'h3a2;
    rom[8566 ] = 12'h3a2;
    rom[8567 ] = 12'h3a2;
    rom[8568 ] = 12'h3a2;
    rom[8569 ] = 12'h3a2;
    rom[8570 ] = 12'h3a2;
    rom[8571 ] = 12'h3a2;
    rom[8572 ] = 12'h3a2;
    rom[8573 ] = 12'h3a2;
    rom[8574 ] = 12'h3a2;
    rom[8575 ] = 12'h3a2;
    rom[8576 ] = 12'h3ca;
    rom[8577 ] = 12'h3ca;
    rom[8578 ] = 12'h3ca;
    rom[8579 ] = 12'h3ca;
    rom[8580 ] = 12'h3ca;
    rom[8581 ] = 12'h3ca;
    rom[8582 ] = 12'h3ca;
    rom[8583 ] = 12'h3ca;
    rom[8584 ] = 12'h3ca;
    rom[8585 ] = 12'h3ca;
    rom[8586 ] = 12'h3ca;
    rom[8587 ] = 12'h3ca;
    rom[8588 ] = 12'h3ca;
    rom[8589 ] = 12'h3ca;
    rom[8590 ] = 12'h3ca;
    rom[8591 ] = 12'h000;
    rom[8592 ] = 12'h000;
    rom[8593 ] = 12'h000;
    rom[8594 ] = 12'h000;
    rom[8595 ] = 12'h000;
    rom[8596 ] = 12'h000;
    rom[8597 ] = 12'h000;
    rom[8598 ] = 12'h000;
    rom[8599 ] = 12'h000;
    rom[8600 ] = 12'h000;
    rom[8601 ] = 12'h000;
    rom[8602 ] = 12'h000;
    rom[8603 ] = 12'h000;
    rom[8604 ] = 12'h000;
    rom[8605 ] = 12'h000;
    rom[8606 ] = 12'h000;
    rom[8607 ] = 12'h000;
    rom[8608 ] = 12'h000;
    rom[8609 ] = 12'h000;
    rom[8610 ] = 12'h000;
    rom[8611 ] = 12'h000;
    rom[8612 ] = 12'h000;
    rom[8613 ] = 12'h000;
    rom[8614 ] = 12'h000;
    rom[8615 ] = 12'h000;
    rom[8616 ] = 12'h000;
    rom[8617 ] = 12'h000;
    rom[8618 ] = 12'h000;
    rom[8619 ] = 12'h3a2;
    rom[8620 ] = 12'h3a2;
    rom[8621 ] = 12'h3a2;
    rom[8622 ] = 12'h3a2;
    rom[8623 ] = 12'h3a2;
    rom[8624 ] = 12'h3a2;
    rom[8625 ] = 12'h3a2;
    rom[8626 ] = 12'h3a2;
    rom[8627 ] = 12'h3a2;
    rom[8628 ] = 12'h3a2;
    rom[8629 ] = 12'h3a2;
    rom[8630 ] = 12'h3a2;
    rom[8631 ] = 12'h3a2;
    rom[8632 ] = 12'h3a2;
    rom[8633 ] = 12'h3a2;
    rom[8634 ] = 12'h3a2;
    rom[8635 ] = 12'h3a2;
    rom[8636 ] = 12'h3a2;
    rom[8637 ] = 12'h3a2;
    rom[8638 ] = 12'h3a2;
    rom[8639 ] = 12'h3a2;
    rom[8640 ] = 12'h3a2;
    rom[8641 ] = 12'h3a2;
    rom[8642 ] = 12'h3a2;
    rom[8643 ] = 12'h3a2;
    rom[8644 ] = 12'h3a2;
    rom[8645 ] = 12'h3a2;
    rom[8646 ] = 12'h3a2;
    rom[8647 ] = 12'h3a2;
    rom[8648 ] = 12'h3a2;
    rom[8649 ] = 12'h3a2;
    rom[8650 ] = 12'h3a2;
    rom[8651 ] = 12'h3a2;
    rom[8652 ] = 12'h3a2;
    rom[8653 ] = 12'h3a2;
    rom[8654 ] = 12'h3a2;
    rom[8655 ] = 12'h3a2;
    rom[8656 ] = 12'h3a2;
    rom[8657 ] = 12'h3a2;
    rom[8658 ] = 12'h000;
    rom[8659 ] = 12'h000;
    rom[8660 ] = 12'h000;
    rom[8661 ] = 12'h000;
    rom[8662 ] = 12'h000;
    rom[8663 ] = 12'h000;
    rom[8664 ] = 12'h000;
    rom[8665 ] = 12'h000;
    rom[8666 ] = 12'h000;
    rom[8667 ] = 12'h000;
    rom[8668 ] = 12'h000;
    rom[8669 ] = 12'h000;
    rom[8670 ] = 12'h000;
    rom[8671 ] = 12'h000;
    rom[8672 ] = 12'h000;
    rom[8673 ] = 12'h000;
    rom[8674 ] = 12'h000;
    rom[8675 ] = 12'h000;
    rom[8676 ] = 12'h000;
    rom[8677 ] = 12'h000;
    rom[8678 ] = 12'h000;
    rom[8679 ] = 12'h000;
    rom[8680 ] = 12'h000;
    rom[8681 ] = 12'h000;
    rom[8682 ] = 12'h000;
    rom[8683 ] = 12'h000;
    rom[8684 ] = 12'h000;
    rom[8685 ] = 12'h000;
    rom[8686 ] = 12'h000;
    rom[8687 ] = 12'h000;
    rom[8688 ] = 12'h000;
    rom[8689 ] = 12'h3a2;
    rom[8690 ] = 12'h3a2;
    rom[8691 ] = 12'h3a2;
    rom[8692 ] = 12'h3a2;
    rom[8693 ] = 12'h3a2;
    rom[8694 ] = 12'h3a2;
    rom[8695 ] = 12'h3a2;
    rom[8696 ] = 12'h3a2;
    rom[8697 ] = 12'h3a2;
    rom[8698 ] = 12'h3a2;
    rom[8699 ] = 12'h3a2;
    rom[8700 ] = 12'h3a2;
    rom[8701 ] = 12'h3a2;
    rom[8702 ] = 12'h3a2;
    rom[8703 ] = 12'h3a2;
    rom[8704 ] = 12'h3ca;
    rom[8705 ] = 12'h3ca;
    rom[8706 ] = 12'h3ca;
    rom[8707 ] = 12'h3ca;
    rom[8708 ] = 12'h3ca;
    rom[8709 ] = 12'h3ca;
    rom[8710 ] = 12'h3ca;
    rom[8711 ] = 12'h3ca;
    rom[8712 ] = 12'h3ca;
    rom[8713 ] = 12'h3ca;
    rom[8714 ] = 12'h3ca;
    rom[8715 ] = 12'h3ca;
    rom[8716 ] = 12'h3da;
    rom[8717 ] = 12'h3da;
    rom[8718 ] = 12'h3da;
    rom[8719 ] = 12'h000;
    rom[8720 ] = 12'h000;
    rom[8721 ] = 12'h000;
    rom[8722 ] = 12'h000;
    rom[8723 ] = 12'h000;
    rom[8724 ] = 12'h000;
    rom[8725 ] = 12'h000;
    rom[8726 ] = 12'h000;
    rom[8727 ] = 12'h000;
    rom[8728 ] = 12'h000;
    rom[8729 ] = 12'h000;
    rom[8730 ] = 12'h000;
    rom[8731 ] = 12'h000;
    rom[8732 ] = 12'h000;
    rom[8733 ] = 12'h000;
    rom[8734 ] = 12'h000;
    rom[8735 ] = 12'h000;
    rom[8736 ] = 12'h000;
    rom[8737 ] = 12'h000;
    rom[8738 ] = 12'h000;
    rom[8739 ] = 12'h000;
    rom[8740 ] = 12'h000;
    rom[8741 ] = 12'h000;
    rom[8742 ] = 12'h000;
    rom[8743 ] = 12'h000;
    rom[8744 ] = 12'h000;
    rom[8745 ] = 12'h000;
    rom[8746 ] = 12'h000;
    rom[8747 ] = 12'h000;
    rom[8748 ] = 12'h391;
    rom[8749 ] = 12'h3a2;
    rom[8750 ] = 12'h3a2;
    rom[8751 ] = 12'h3a2;
    rom[8752 ] = 12'h3a2;
    rom[8753 ] = 12'h3a2;
    rom[8754 ] = 12'h3a2;
    rom[8755 ] = 12'h3a2;
    rom[8756 ] = 12'h3a2;
    rom[8757 ] = 12'h3a2;
    rom[8758 ] = 12'h3a2;
    rom[8759 ] = 12'h3a2;
    rom[8760 ] = 12'h3a2;
    rom[8761 ] = 12'h3a2;
    rom[8762 ] = 12'h3a2;
    rom[8763 ] = 12'h3a2;
    rom[8764 ] = 12'h3a2;
    rom[8765 ] = 12'h3a2;
    rom[8766 ] = 12'h3a2;
    rom[8767 ] = 12'h3a2;
    rom[8768 ] = 12'h3a2;
    rom[8769 ] = 12'h3a2;
    rom[8770 ] = 12'h3a2;
    rom[8771 ] = 12'h3a2;
    rom[8772 ] = 12'h3a2;
    rom[8773 ] = 12'h3a2;
    rom[8774 ] = 12'h3a2;
    rom[8775 ] = 12'h3a2;
    rom[8776 ] = 12'h3a2;
    rom[8777 ] = 12'h3a2;
    rom[8778 ] = 12'h3a2;
    rom[8779 ] = 12'h3a2;
    rom[8780 ] = 12'h3a2;
    rom[8781 ] = 12'h3a2;
    rom[8782 ] = 12'h3a2;
    rom[8783 ] = 12'h3a2;
    rom[8784 ] = 12'h392;
    rom[8785 ] = 12'h000;
    rom[8786 ] = 12'h000;
    rom[8787 ] = 12'h000;
    rom[8788 ] = 12'h000;
    rom[8789 ] = 12'h000;
    rom[8790 ] = 12'h000;
    rom[8791 ] = 12'h000;
    rom[8792 ] = 12'h000;
    rom[8793 ] = 12'h000;
    rom[8794 ] = 12'h000;
    rom[8795 ] = 12'h000;
    rom[8796 ] = 12'h000;
    rom[8797 ] = 12'h000;
    rom[8798 ] = 12'h000;
    rom[8799 ] = 12'h000;
    rom[8800 ] = 12'h000;
    rom[8801 ] = 12'h000;
    rom[8802 ] = 12'h000;
    rom[8803 ] = 12'h000;
    rom[8804 ] = 12'h000;
    rom[8805 ] = 12'h000;
    rom[8806 ] = 12'h000;
    rom[8807 ] = 12'h000;
    rom[8808 ] = 12'h000;
    rom[8809 ] = 12'h000;
    rom[8810 ] = 12'h000;
    rom[8811 ] = 12'h000;
    rom[8812 ] = 12'h000;
    rom[8813 ] = 12'h000;
    rom[8814 ] = 12'h000;
    rom[8815 ] = 12'h000;
    rom[8816 ] = 12'h000;
    rom[8817 ] = 12'h3a2;
    rom[8818 ] = 12'h3a2;
    rom[8819 ] = 12'h3a2;
    rom[8820 ] = 12'h3a2;
    rom[8821 ] = 12'h3a2;
    rom[8822 ] = 12'h3a2;
    rom[8823 ] = 12'h3a2;
    rom[8824 ] = 12'h3a2;
    rom[8825 ] = 12'h3a2;
    rom[8826 ] = 12'h3a2;
    rom[8827 ] = 12'h3a2;
    rom[8828 ] = 12'h3a2;
    rom[8829 ] = 12'h3a2;
    rom[8830 ] = 12'h3a2;
    rom[8831 ] = 12'h3a2;
    rom[8832 ] = 12'h3ca;
    rom[8833 ] = 12'h3ca;
    rom[8834 ] = 12'h3ca;
    rom[8835 ] = 12'h3ca;
    rom[8836 ] = 12'h3ca;
    rom[8837 ] = 12'h3ca;
    rom[8838 ] = 12'h3ca;
    rom[8839 ] = 12'h3ca;
    rom[8840 ] = 12'h3ca;
    rom[8841 ] = 12'h3da;
    rom[8842 ] = 12'h3da;
    rom[8843 ] = 12'h3da;
    rom[8844 ] = 12'h3da;
    rom[8845 ] = 12'h3da;
    rom[8846 ] = 12'h3da;
    rom[8847 ] = 12'h000;
    rom[8848 ] = 12'h000;
    rom[8849 ] = 12'h000;
    rom[8850 ] = 12'h000;
    rom[8851 ] = 12'h000;
    rom[8852 ] = 12'h000;
    rom[8853 ] = 12'h000;
    rom[8854 ] = 12'h000;
    rom[8855 ] = 12'h000;
    rom[8856 ] = 12'h000;
    rom[8857 ] = 12'h000;
    rom[8858 ] = 12'h000;
    rom[8859 ] = 12'h000;
    rom[8860 ] = 12'h000;
    rom[8861 ] = 12'h000;
    rom[8862 ] = 12'h000;
    rom[8863 ] = 12'h000;
    rom[8864 ] = 12'h000;
    rom[8865 ] = 12'h000;
    rom[8866 ] = 12'h000;
    rom[8867 ] = 12'h000;
    rom[8868 ] = 12'h000;
    rom[8869 ] = 12'h000;
    rom[8870 ] = 12'h000;
    rom[8871 ] = 12'h000;
    rom[8872 ] = 12'h000;
    rom[8873 ] = 12'h000;
    rom[8874 ] = 12'h000;
    rom[8875 ] = 12'h000;
    rom[8876 ] = 12'h000;
    rom[8877 ] = 12'h000;
    rom[8878 ] = 12'h3a2;
    rom[8879 ] = 12'h3a2;
    rom[8880 ] = 12'h3a2;
    rom[8881 ] = 12'h3a2;
    rom[8882 ] = 12'h3a2;
    rom[8883 ] = 12'h3a2;
    rom[8884 ] = 12'h3a2;
    rom[8885 ] = 12'h3a2;
    rom[8886 ] = 12'h3a2;
    rom[8887 ] = 12'h3a2;
    rom[8888 ] = 12'h3a2;
    rom[8889 ] = 12'h3a2;
    rom[8890 ] = 12'h3a2;
    rom[8891 ] = 12'h3a2;
    rom[8892 ] = 12'h3a2;
    rom[8893 ] = 12'h3a2;
    rom[8894 ] = 12'h3a2;
    rom[8895 ] = 12'h3a2;
    rom[8896 ] = 12'h3a2;
    rom[8897 ] = 12'h3a2;
    rom[8898 ] = 12'h3a2;
    rom[8899 ] = 12'h3a2;
    rom[8900 ] = 12'h3a2;
    rom[8901 ] = 12'h3a2;
    rom[8902 ] = 12'h3a2;
    rom[8903 ] = 12'h3a2;
    rom[8904 ] = 12'h3a2;
    rom[8905 ] = 12'h3a2;
    rom[8906 ] = 12'h3a2;
    rom[8907 ] = 12'h3a2;
    rom[8908 ] = 12'h3a2;
    rom[8909 ] = 12'h3a2;
    rom[8910 ] = 12'h3a2;
    rom[8911 ] = 12'h000;
    rom[8912 ] = 12'h000;
    rom[8913 ] = 12'h000;
    rom[8914 ] = 12'h000;
    rom[8915 ] = 12'h000;
    rom[8916 ] = 12'h000;
    rom[8917 ] = 12'h000;
    rom[8918 ] = 12'h000;
    rom[8919 ] = 12'h000;
    rom[8920 ] = 12'h000;
    rom[8921 ] = 12'h000;
    rom[8922 ] = 12'h000;
    rom[8923 ] = 12'h000;
    rom[8924 ] = 12'h000;
    rom[8925 ] = 12'h000;
    rom[8926 ] = 12'h000;
    rom[8927 ] = 12'h000;
    rom[8928 ] = 12'h000;
    rom[8929 ] = 12'h000;
    rom[8930 ] = 12'h000;
    rom[8931 ] = 12'h000;
    rom[8932 ] = 12'h000;
    rom[8933 ] = 12'h000;
    rom[8934 ] = 12'h000;
    rom[8935 ] = 12'h000;
    rom[8936 ] = 12'h000;
    rom[8937 ] = 12'h000;
    rom[8938 ] = 12'h000;
    rom[8939 ] = 12'h000;
    rom[8940 ] = 12'h000;
    rom[8941 ] = 12'h000;
    rom[8942 ] = 12'h000;
    rom[8943 ] = 12'h000;
    rom[8944 ] = 12'h000;
    rom[8945 ] = 12'h3a2;
    rom[8946 ] = 12'h3a2;
    rom[8947 ] = 12'h3a2;
    rom[8948 ] = 12'h3a2;
    rom[8949 ] = 12'h3a2;
    rom[8950 ] = 12'h3a2;
    rom[8951 ] = 12'h3a2;
    rom[8952 ] = 12'h3a2;
    rom[8953 ] = 12'h3a2;
    rom[8954 ] = 12'h3a2;
    rom[8955 ] = 12'h3a2;
    rom[8956 ] = 12'h3a2;
    rom[8957 ] = 12'h3a2;
    rom[8958 ] = 12'h3a2;
    rom[8959 ] = 12'h3a2;
    rom[8960 ] = 12'h3ca;
    rom[8961 ] = 12'h3ca;
    rom[8962 ] = 12'h3ca;
    rom[8963 ] = 12'h3ca;
    rom[8964 ] = 12'h3ca;
    rom[8965 ] = 12'h3ca;
    rom[8966 ] = 12'h3da;
    rom[8967 ] = 12'h3da;
    rom[8968 ] = 12'h3da;
    rom[8969 ] = 12'h3da;
    rom[8970 ] = 12'h3da;
    rom[8971 ] = 12'h3da;
    rom[8972 ] = 12'h3da;
    rom[8973 ] = 12'h3db;
    rom[8974 ] = 12'h3db;
    rom[8975 ] = 12'h000;
    rom[8976 ] = 12'h000;
    rom[8977 ] = 12'h000;
    rom[8978 ] = 12'h000;
    rom[8979 ] = 12'h000;
    rom[8980 ] = 12'h000;
    rom[8981 ] = 12'h000;
    rom[8982 ] = 12'h000;
    rom[8983 ] = 12'h000;
    rom[8984 ] = 12'h000;
    rom[8985 ] = 12'h000;
    rom[8986 ] = 12'h000;
    rom[8987 ] = 12'h000;
    rom[8988 ] = 12'h000;
    rom[8989 ] = 12'h000;
    rom[8990 ] = 12'h000;
    rom[8991 ] = 12'h000;
    rom[8992 ] = 12'h000;
    rom[8993 ] = 12'h000;
    rom[8994 ] = 12'h000;
    rom[8995 ] = 12'h000;
    rom[8996 ] = 12'h000;
    rom[8997 ] = 12'h000;
    rom[8998 ] = 12'h000;
    rom[8999 ] = 12'h000;
    rom[9000 ] = 12'h000;
    rom[9001 ] = 12'h000;
    rom[9002 ] = 12'h000;
    rom[9003 ] = 12'h000;
    rom[9004 ] = 12'h000;
    rom[9005 ] = 12'h000;
    rom[9006 ] = 12'h000;
    rom[9007 ] = 12'h000;
    rom[9008 ] = 12'h3a2;
    rom[9009 ] = 12'h3a2;
    rom[9010 ] = 12'h3a2;
    rom[9011 ] = 12'h3a2;
    rom[9012 ] = 12'h3a2;
    rom[9013 ] = 12'h3a2;
    rom[9014 ] = 12'h3a2;
    rom[9015 ] = 12'h3a2;
    rom[9016 ] = 12'h3a2;
    rom[9017 ] = 12'h3a2;
    rom[9018 ] = 12'h3a2;
    rom[9019 ] = 12'h3a2;
    rom[9020 ] = 12'h3a2;
    rom[9021 ] = 12'h3a2;
    rom[9022 ] = 12'h3a2;
    rom[9023 ] = 12'h3a2;
    rom[9024 ] = 12'h3a2;
    rom[9025 ] = 12'h3a2;
    rom[9026 ] = 12'h3a2;
    rom[9027 ] = 12'h3a2;
    rom[9028 ] = 12'h3a2;
    rom[9029 ] = 12'h3a2;
    rom[9030 ] = 12'h3a2;
    rom[9031 ] = 12'h3a2;
    rom[9032 ] = 12'h3a2;
    rom[9033 ] = 12'h3a2;
    rom[9034 ] = 12'h3a2;
    rom[9035 ] = 12'h3a2;
    rom[9036 ] = 12'h3a2;
    rom[9037 ] = 12'h3a2;
    rom[9038 ] = 12'h000;
    rom[9039 ] = 12'h000;
    rom[9040 ] = 12'h000;
    rom[9041 ] = 12'h000;
    rom[9042 ] = 12'h000;
    rom[9043 ] = 12'h000;
    rom[9044 ] = 12'h000;
    rom[9045 ] = 12'h000;
    rom[9046 ] = 12'h000;
    rom[9047 ] = 12'h000;
    rom[9048 ] = 12'h000;
    rom[9049 ] = 12'h000;
    rom[9050 ] = 12'h000;
    rom[9051 ] = 12'h000;
    rom[9052 ] = 12'h000;
    rom[9053 ] = 12'h000;
    rom[9054 ] = 12'h000;
    rom[9055 ] = 12'h000;
    rom[9056 ] = 12'h000;
    rom[9057 ] = 12'h000;
    rom[9058 ] = 12'h000;
    rom[9059 ] = 12'h000;
    rom[9060 ] = 12'h000;
    rom[9061 ] = 12'h000;
    rom[9062 ] = 12'h000;
    rom[9063 ] = 12'h000;
    rom[9064 ] = 12'h000;
    rom[9065 ] = 12'h000;
    rom[9066 ] = 12'h000;
    rom[9067 ] = 12'h000;
    rom[9068 ] = 12'h000;
    rom[9069 ] = 12'h000;
    rom[9070 ] = 12'h000;
    rom[9071 ] = 12'h000;
    rom[9072 ] = 12'h000;
    rom[9073 ] = 12'h3a2;
    rom[9074 ] = 12'h3a2;
    rom[9075 ] = 12'h3a2;
    rom[9076 ] = 12'h3a2;
    rom[9077 ] = 12'h3a2;
    rom[9078 ] = 12'h3a2;
    rom[9079 ] = 12'h3a2;
    rom[9080 ] = 12'h3a2;
    rom[9081 ] = 12'h3a2;
    rom[9082 ] = 12'h3a2;
    rom[9083 ] = 12'h3a2;
    rom[9084 ] = 12'h3a2;
    rom[9085 ] = 12'h3a2;
    rom[9086 ] = 12'h3a2;
    rom[9087 ] = 12'h3a2;
    rom[9088 ] = 12'h3ca;
    rom[9089 ] = 12'h3ca;
    rom[9090 ] = 12'h3ca;
    rom[9091 ] = 12'h3da;
    rom[9092 ] = 12'h3da;
    rom[9093 ] = 12'h3da;
    rom[9094 ] = 12'h3da;
    rom[9095 ] = 12'h3da;
    rom[9096 ] = 12'h3da;
    rom[9097 ] = 12'h3da;
    rom[9098 ] = 12'h3db;
    rom[9099 ] = 12'h3db;
    rom[9100 ] = 12'h3db;
    rom[9101 ] = 12'h3db;
    rom[9102 ] = 12'h3db;
    rom[9103 ] = 12'h000;
    rom[9104 ] = 12'h000;
    rom[9105 ] = 12'h000;
    rom[9106 ] = 12'h000;
    rom[9107 ] = 12'h000;
    rom[9108 ] = 12'h000;
    rom[9109 ] = 12'h000;
    rom[9110 ] = 12'h000;
    rom[9111 ] = 12'h000;
    rom[9112 ] = 12'h000;
    rom[9113 ] = 12'h000;
    rom[9114 ] = 12'h000;
    rom[9115 ] = 12'h000;
    rom[9116 ] = 12'h000;
    rom[9117 ] = 12'h000;
    rom[9118 ] = 12'h000;
    rom[9119 ] = 12'h000;
    rom[9120 ] = 12'h000;
    rom[9121 ] = 12'h000;
    rom[9122 ] = 12'h000;
    rom[9123 ] = 12'h000;
    rom[9124 ] = 12'h000;
    rom[9125 ] = 12'h000;
    rom[9126 ] = 12'h000;
    rom[9127 ] = 12'h000;
    rom[9128 ] = 12'h000;
    rom[9129 ] = 12'h000;
    rom[9130 ] = 12'h000;
    rom[9131 ] = 12'h000;
    rom[9132 ] = 12'h000;
    rom[9133 ] = 12'h000;
    rom[9134 ] = 12'h000;
    rom[9135 ] = 12'h000;
    rom[9136 ] = 12'h000;
    rom[9137 ] = 12'h3a2;
    rom[9138 ] = 12'h3a2;
    rom[9139 ] = 12'h3a2;
    rom[9140 ] = 12'h3a2;
    rom[9141 ] = 12'h3a2;
    rom[9142 ] = 12'h3a2;
    rom[9143 ] = 12'h3a2;
    rom[9144 ] = 12'h3a2;
    rom[9145 ] = 12'h3a2;
    rom[9146 ] = 12'h3a2;
    rom[9147 ] = 12'h3a2;
    rom[9148 ] = 12'h3a2;
    rom[9149 ] = 12'h3a2;
    rom[9150 ] = 12'h3a2;
    rom[9151 ] = 12'h3a2;
    rom[9152 ] = 12'h3a2;
    rom[9153 ] = 12'h3a2;
    rom[9154 ] = 12'h3a2;
    rom[9155 ] = 12'h3a2;
    rom[9156 ] = 12'h3a2;
    rom[9157 ] = 12'h3a2;
    rom[9158 ] = 12'h3a2;
    rom[9159 ] = 12'h3a2;
    rom[9160 ] = 12'h3a2;
    rom[9161 ] = 12'h3a2;
    rom[9162 ] = 12'h3a2;
    rom[9163 ] = 12'h3a2;
    rom[9164 ] = 12'h3a2;
    rom[9165 ] = 12'h000;
    rom[9166 ] = 12'h000;
    rom[9167 ] = 12'h000;
    rom[9168 ] = 12'h000;
    rom[9169 ] = 12'h000;
    rom[9170 ] = 12'h000;
    rom[9171 ] = 12'h000;
    rom[9172 ] = 12'h000;
    rom[9173 ] = 12'h000;
    rom[9174 ] = 12'h000;
    rom[9175 ] = 12'h000;
    rom[9176 ] = 12'h000;
    rom[9177 ] = 12'h000;
    rom[9178 ] = 12'h000;
    rom[9179 ] = 12'h000;
    rom[9180 ] = 12'h000;
    rom[9181 ] = 12'h000;
    rom[9182 ] = 12'h000;
    rom[9183 ] = 12'h000;
    rom[9184 ] = 12'h000;
    rom[9185 ] = 12'h000;
    rom[9186 ] = 12'h000;
    rom[9187 ] = 12'h000;
    rom[9188 ] = 12'h000;
    rom[9189 ] = 12'h000;
    rom[9190 ] = 12'h000;
    rom[9191 ] = 12'h000;
    rom[9192 ] = 12'h000;
    rom[9193 ] = 12'h000;
    rom[9194 ] = 12'h000;
    rom[9195 ] = 12'h000;
    rom[9196 ] = 12'h000;
    rom[9197 ] = 12'h000;
    rom[9198 ] = 12'h000;
    rom[9199 ] = 12'h000;
    rom[9200 ] = 12'h000;
    rom[9201 ] = 12'h3a2;
    rom[9202 ] = 12'h3a2;
    rom[9203 ] = 12'h3a2;
    rom[9204 ] = 12'h3a2;
    rom[9205 ] = 12'h3a2;
    rom[9206 ] = 12'h3a2;
    rom[9207 ] = 12'h3a2;
    rom[9208 ] = 12'h3a2;
    rom[9209 ] = 12'h3a2;
    rom[9210 ] = 12'h3a2;
    rom[9211 ] = 12'h3a2;
    rom[9212 ] = 12'h3a2;
    rom[9213 ] = 12'h3a2;
    rom[9214 ] = 12'h3a2;
    rom[9215 ] = 12'h3a2;
    rom[9216 ] = 12'h3c9;
    rom[9217 ] = 12'h3da;
    rom[9218 ] = 12'h3da;
    rom[9219 ] = 12'h3da;
    rom[9220 ] = 12'h3da;
    rom[9221 ] = 12'h3da;
    rom[9222 ] = 12'h3da;
    rom[9223 ] = 12'h3db;
    rom[9224 ] = 12'h3db;
    rom[9225 ] = 12'h3db;
    rom[9226 ] = 12'h3db;
    rom[9227 ] = 12'h3db;
    rom[9228 ] = 12'h3db;
    rom[9229 ] = 12'h3db;
    rom[9230 ] = 12'h3db;
    rom[9231 ] = 12'h2db;
    rom[9232 ] = 12'h000;
    rom[9233 ] = 12'h000;
    rom[9234 ] = 12'h000;
    rom[9235 ] = 12'h000;
    rom[9236 ] = 12'h000;
    rom[9237 ] = 12'h000;
    rom[9238 ] = 12'h000;
    rom[9239 ] = 12'h000;
    rom[9240 ] = 12'h000;
    rom[9241 ] = 12'h000;
    rom[9242 ] = 12'h000;
    rom[9243 ] = 12'h000;
    rom[9244 ] = 12'h000;
    rom[9245 ] = 12'h000;
    rom[9246 ] = 12'h000;
    rom[9247 ] = 12'h000;
    rom[9248 ] = 12'h000;
    rom[9249 ] = 12'h000;
    rom[9250 ] = 12'h000;
    rom[9251 ] = 12'h000;
    rom[9252 ] = 12'h000;
    rom[9253 ] = 12'h000;
    rom[9254 ] = 12'h000;
    rom[9255 ] = 12'h000;
    rom[9256 ] = 12'h000;
    rom[9257 ] = 12'h000;
    rom[9258 ] = 12'h000;
    rom[9259 ] = 12'h000;
    rom[9260 ] = 12'h000;
    rom[9261 ] = 12'h000;
    rom[9262 ] = 12'h000;
    rom[9263 ] = 12'h000;
    rom[9264 ] = 12'h000;
    rom[9265 ] = 12'h000;
    rom[9266 ] = 12'h000;
    rom[9267 ] = 12'h3a2;
    rom[9268 ] = 12'h3a2;
    rom[9269 ] = 12'h3a2;
    rom[9270 ] = 12'h3a2;
    rom[9271 ] = 12'h3a2;
    rom[9272 ] = 12'h3a2;
    rom[9273 ] = 12'h3a2;
    rom[9274 ] = 12'h3a2;
    rom[9275 ] = 12'h3a2;
    rom[9276 ] = 12'h3a2;
    rom[9277 ] = 12'h3a2;
    rom[9278 ] = 12'h3a2;
    rom[9279 ] = 12'h3a2;
    rom[9280 ] = 12'h3a2;
    rom[9281 ] = 12'h3a2;
    rom[9282 ] = 12'h3a2;
    rom[9283 ] = 12'h3a2;
    rom[9284 ] = 12'h3a2;
    rom[9285 ] = 12'h3a2;
    rom[9286 ] = 12'h3a2;
    rom[9287 ] = 12'h3a2;
    rom[9288 ] = 12'h3a2;
    rom[9289 ] = 12'h3a2;
    rom[9290 ] = 12'h3a2;
    rom[9291 ] = 12'h000;
    rom[9292 ] = 12'h000;
    rom[9293 ] = 12'h000;
    rom[9294 ] = 12'h000;
    rom[9295 ] = 12'h000;
    rom[9296 ] = 12'h000;
    rom[9297 ] = 12'h000;
    rom[9298 ] = 12'h000;
    rom[9299 ] = 12'h000;
    rom[9300 ] = 12'h000;
    rom[9301 ] = 12'h000;
    rom[9302 ] = 12'h000;
    rom[9303 ] = 12'h000;
    rom[9304 ] = 12'h000;
    rom[9305 ] = 12'h000;
    rom[9306 ] = 12'h000;
    rom[9307 ] = 12'h000;
    rom[9308 ] = 12'h000;
    rom[9309 ] = 12'h000;
    rom[9310 ] = 12'h000;
    rom[9311 ] = 12'h000;
    rom[9312 ] = 12'h000;
    rom[9313 ] = 12'h000;
    rom[9314 ] = 12'h000;
    rom[9315 ] = 12'h000;
    rom[9316 ] = 12'h000;
    rom[9317 ] = 12'h000;
    rom[9318 ] = 12'h000;
    rom[9319 ] = 12'h000;
    rom[9320 ] = 12'h000;
    rom[9321 ] = 12'h000;
    rom[9322 ] = 12'h000;
    rom[9323 ] = 12'h000;
    rom[9324 ] = 12'h000;
    rom[9325 ] = 12'h000;
    rom[9326 ] = 12'h000;
    rom[9327 ] = 12'h000;
    rom[9328 ] = 12'h3a2;
    rom[9329 ] = 12'h3a2;
    rom[9330 ] = 12'h3a2;
    rom[9331 ] = 12'h3a2;
    rom[9332 ] = 12'h3a2;
    rom[9333 ] = 12'h3a2;
    rom[9334 ] = 12'h3a2;
    rom[9335 ] = 12'h3a2;
    rom[9336 ] = 12'h3a2;
    rom[9337 ] = 12'h3a2;
    rom[9338 ] = 12'h3a2;
    rom[9339 ] = 12'h3a2;
    rom[9340 ] = 12'h3a2;
    rom[9341 ] = 12'h3a2;
    rom[9342 ] = 12'h3a2;
    rom[9343 ] = 12'h3a2;
    rom[9344 ] = 12'h000;
    rom[9345 ] = 12'h3da;
    rom[9346 ] = 12'h3da;
    rom[9347 ] = 12'h3da;
    rom[9348 ] = 12'h3db;
    rom[9349 ] = 12'h3db;
    rom[9350 ] = 12'h3db;
    rom[9351 ] = 12'h3db;
    rom[9352 ] = 12'h3db;
    rom[9353 ] = 12'h3db;
    rom[9354 ] = 12'h3db;
    rom[9355 ] = 12'h3db;
    rom[9356 ] = 12'h2db;
    rom[9357 ] = 12'h2db;
    rom[9358 ] = 12'h2db;
    rom[9359 ] = 12'h2db;
    rom[9360 ] = 12'h000;
    rom[9361 ] = 12'h000;
    rom[9362 ] = 12'h000;
    rom[9363 ] = 12'h000;
    rom[9364 ] = 12'h000;
    rom[9365 ] = 12'h000;
    rom[9366 ] = 12'h000;
    rom[9367 ] = 12'h000;
    rom[9368 ] = 12'h000;
    rom[9369 ] = 12'h000;
    rom[9370 ] = 12'h000;
    rom[9371 ] = 12'h000;
    rom[9372 ] = 12'h000;
    rom[9373 ] = 12'h000;
    rom[9374 ] = 12'h000;
    rom[9375 ] = 12'h000;
    rom[9376 ] = 12'h000;
    rom[9377 ] = 12'h000;
    rom[9378 ] = 12'h000;
    rom[9379 ] = 12'h000;
    rom[9380 ] = 12'h000;
    rom[9381 ] = 12'h000;
    rom[9382 ] = 12'h000;
    rom[9383 ] = 12'h000;
    rom[9384 ] = 12'h000;
    rom[9385 ] = 12'h000;
    rom[9386 ] = 12'h000;
    rom[9387 ] = 12'h000;
    rom[9388 ] = 12'h000;
    rom[9389 ] = 12'h000;
    rom[9390 ] = 12'h000;
    rom[9391 ] = 12'h000;
    rom[9392 ] = 12'h000;
    rom[9393 ] = 12'h000;
    rom[9394 ] = 12'h000;
    rom[9395 ] = 12'h000;
    rom[9396 ] = 12'h392;
    rom[9397 ] = 12'h3a2;
    rom[9398 ] = 12'h3a2;
    rom[9399 ] = 12'h3a2;
    rom[9400 ] = 12'h3a2;
    rom[9401 ] = 12'h3a2;
    rom[9402 ] = 12'h3a2;
    rom[9403 ] = 12'h3a2;
    rom[9404 ] = 12'h3a2;
    rom[9405 ] = 12'h3a2;
    rom[9406 ] = 12'h3a2;
    rom[9407 ] = 12'h3a2;
    rom[9408 ] = 12'h3a2;
    rom[9409 ] = 12'h3a2;
    rom[9410 ] = 12'h3a2;
    rom[9411 ] = 12'h3a2;
    rom[9412 ] = 12'h3a2;
    rom[9413 ] = 12'h3a2;
    rom[9414 ] = 12'h3a2;
    rom[9415 ] = 12'h3a2;
    rom[9416 ] = 12'h3a2;
    rom[9417 ] = 12'h3a2;
    rom[9418 ] = 12'h000;
    rom[9419 ] = 12'h000;
    rom[9420 ] = 12'h000;
    rom[9421 ] = 12'h000;
    rom[9422 ] = 12'h000;
    rom[9423 ] = 12'h000;
    rom[9424 ] = 12'h000;
    rom[9425 ] = 12'h000;
    rom[9426 ] = 12'h000;
    rom[9427 ] = 12'h000;
    rom[9428 ] = 12'h000;
    rom[9429 ] = 12'h000;
    rom[9430 ] = 12'h000;
    rom[9431 ] = 12'h000;
    rom[9432 ] = 12'h000;
    rom[9433 ] = 12'h000;
    rom[9434 ] = 12'h000;
    rom[9435 ] = 12'h000;
    rom[9436 ] = 12'h000;
    rom[9437 ] = 12'h000;
    rom[9438 ] = 12'h000;
    rom[9439 ] = 12'h000;
    rom[9440 ] = 12'h000;
    rom[9441 ] = 12'h000;
    rom[9442 ] = 12'h000;
    rom[9443 ] = 12'h000;
    rom[9444 ] = 12'h000;
    rom[9445 ] = 12'h000;
    rom[9446 ] = 12'h000;
    rom[9447 ] = 12'h000;
    rom[9448 ] = 12'h000;
    rom[9449 ] = 12'h000;
    rom[9450 ] = 12'h000;
    rom[9451 ] = 12'h000;
    rom[9452 ] = 12'h000;
    rom[9453 ] = 12'h000;
    rom[9454 ] = 12'h000;
    rom[9455 ] = 12'h000;
    rom[9456 ] = 12'h3a2;
    rom[9457 ] = 12'h3a2;
    rom[9458 ] = 12'h3a2;
    rom[9459 ] = 12'h3a2;
    rom[9460 ] = 12'h3a2;
    rom[9461 ] = 12'h3a2;
    rom[9462 ] = 12'h3a2;
    rom[9463 ] = 12'h3a2;
    rom[9464 ] = 12'h3a2;
    rom[9465 ] = 12'h3a2;
    rom[9466 ] = 12'h3a2;
    rom[9467 ] = 12'h3a2;
    rom[9468 ] = 12'h3a2;
    rom[9469 ] = 12'h3a2;
    rom[9470 ] = 12'h3a2;
    rom[9471 ] = 12'h000;
    rom[9472 ] = 12'h000;
    rom[9473 ] = 12'h3db;
    rom[9474 ] = 12'h3db;
    rom[9475 ] = 12'h3db;
    rom[9476 ] = 12'h3db;
    rom[9477 ] = 12'h3db;
    rom[9478 ] = 12'h3db;
    rom[9479 ] = 12'h3db;
    rom[9480 ] = 12'h3db;
    rom[9481 ] = 12'h2db;
    rom[9482 ] = 12'h2db;
    rom[9483 ] = 12'h2db;
    rom[9484 ] = 12'h2db;
    rom[9485 ] = 12'h2db;
    rom[9486 ] = 12'h2db;
    rom[9487 ] = 12'h2db;
    rom[9488 ] = 12'h000;
    rom[9489 ] = 12'h000;
    rom[9490 ] = 12'h000;
    rom[9491 ] = 12'h000;
    rom[9492 ] = 12'h000;
    rom[9493 ] = 12'h000;
    rom[9494 ] = 12'h000;
    rom[9495 ] = 12'h000;
    rom[9496 ] = 12'h000;
    rom[9497 ] = 12'h000;
    rom[9498 ] = 12'h000;
    rom[9499 ] = 12'h000;
    rom[9500 ] = 12'h000;
    rom[9501 ] = 12'h000;
    rom[9502 ] = 12'h000;
    rom[9503 ] = 12'h000;
    rom[9504 ] = 12'h000;
    rom[9505 ] = 12'h000;
    rom[9506 ] = 12'h000;
    rom[9507 ] = 12'h000;
    rom[9508 ] = 12'h000;
    rom[9509 ] = 12'h000;
    rom[9510 ] = 12'h000;
    rom[9511 ] = 12'h000;
    rom[9512 ] = 12'h000;
    rom[9513 ] = 12'h000;
    rom[9514 ] = 12'h000;
    rom[9515 ] = 12'h000;
    rom[9516 ] = 12'h000;
    rom[9517 ] = 12'h000;
    rom[9518 ] = 12'h000;
    rom[9519 ] = 12'h000;
    rom[9520 ] = 12'h000;
    rom[9521 ] = 12'h000;
    rom[9522 ] = 12'h000;
    rom[9523 ] = 12'h000;
    rom[9524 ] = 12'h000;
    rom[9525 ] = 12'h000;
    rom[9526 ] = 12'h3a2;
    rom[9527 ] = 12'h3a2;
    rom[9528 ] = 12'h3a2;
    rom[9529 ] = 12'h3a2;
    rom[9530 ] = 12'h3a2;
    rom[9531 ] = 12'h3a2;
    rom[9532 ] = 12'h3a2;
    rom[9533 ] = 12'h3a2;
    rom[9534 ] = 12'h3a2;
    rom[9535 ] = 12'h3a2;
    rom[9536 ] = 12'h3a2;
    rom[9537 ] = 12'h3a2;
    rom[9538 ] = 12'h3a2;
    rom[9539 ] = 12'h3a2;
    rom[9540 ] = 12'h3a2;
    rom[9541 ] = 12'h3a2;
    rom[9542 ] = 12'h3a2;
    rom[9543 ] = 12'h3a2;
    rom[9544 ] = 12'h3a2;
    rom[9545 ] = 12'h000;
    rom[9546 ] = 12'h000;
    rom[9547 ] = 12'h000;
    rom[9548 ] = 12'h000;
    rom[9549 ] = 12'h000;
    rom[9550 ] = 12'h000;
    rom[9551 ] = 12'h000;
    rom[9552 ] = 12'h000;
    rom[9553 ] = 12'h000;
    rom[9554 ] = 12'h000;
    rom[9555 ] = 12'h000;
    rom[9556 ] = 12'h000;
    rom[9557 ] = 12'h000;
    rom[9558 ] = 12'h000;
    rom[9559 ] = 12'h000;
    rom[9560 ] = 12'h000;
    rom[9561 ] = 12'h000;
    rom[9562 ] = 12'h000;
    rom[9563 ] = 12'h000;
    rom[9564 ] = 12'h000;
    rom[9565 ] = 12'h000;
    rom[9566 ] = 12'h000;
    rom[9567 ] = 12'h000;
    rom[9568 ] = 12'h000;
    rom[9569 ] = 12'h000;
    rom[9570 ] = 12'h000;
    rom[9571 ] = 12'h000;
    rom[9572 ] = 12'h000;
    rom[9573 ] = 12'h000;
    rom[9574 ] = 12'h000;
    rom[9575 ] = 12'h000;
    rom[9576 ] = 12'h000;
    rom[9577 ] = 12'h000;
    rom[9578 ] = 12'h000;
    rom[9579 ] = 12'h000;
    rom[9580 ] = 12'h000;
    rom[9581 ] = 12'h000;
    rom[9582 ] = 12'h000;
    rom[9583 ] = 12'h000;
    rom[9584 ] = 12'h3a2;
    rom[9585 ] = 12'h3a2;
    rom[9586 ] = 12'h3a2;
    rom[9587 ] = 12'h3a2;
    rom[9588 ] = 12'h3a2;
    rom[9589 ] = 12'h3a2;
    rom[9590 ] = 12'h3a2;
    rom[9591 ] = 12'h3a2;
    rom[9592 ] = 12'h3a2;
    rom[9593 ] = 12'h3a2;
    rom[9594 ] = 12'h3a2;
    rom[9595 ] = 12'h3a2;
    rom[9596 ] = 12'h3a2;
    rom[9597 ] = 12'h3a2;
    rom[9598 ] = 12'h3a2;
    rom[9599 ] = 12'h000;
    rom[9600 ] = 12'h000;
    rom[9601 ] = 12'h3db;
    rom[9602 ] = 12'h3db;
    rom[9603 ] = 12'h3db;
    rom[9604 ] = 12'h3db;
    rom[9605 ] = 12'h3db;
    rom[9606 ] = 12'h2db;
    rom[9607 ] = 12'h2db;
    rom[9608 ] = 12'h2db;
    rom[9609 ] = 12'h2db;
    rom[9610 ] = 12'h2db;
    rom[9611 ] = 12'h2db;
    rom[9612 ] = 12'h2db;
    rom[9613 ] = 12'h2db;
    rom[9614 ] = 12'h2db;
    rom[9615 ] = 12'h2db;
    rom[9616 ] = 12'h000;
    rom[9617 ] = 12'h000;
    rom[9618 ] = 12'h000;
    rom[9619 ] = 12'h000;
    rom[9620 ] = 12'h000;
    rom[9621 ] = 12'h000;
    rom[9622 ] = 12'h000;
    rom[9623 ] = 12'h000;
    rom[9624 ] = 12'h000;
    rom[9625 ] = 12'h000;
    rom[9626 ] = 12'h000;
    rom[9627 ] = 12'h000;
    rom[9628 ] = 12'h000;
    rom[9629 ] = 12'h000;
    rom[9630 ] = 12'h000;
    rom[9631 ] = 12'h000;
    rom[9632 ] = 12'h000;
    rom[9633 ] = 12'h000;
    rom[9634 ] = 12'h000;
    rom[9635 ] = 12'h000;
    rom[9636 ] = 12'h000;
    rom[9637 ] = 12'h000;
    rom[9638 ] = 12'h000;
    rom[9639 ] = 12'h000;
    rom[9640 ] = 12'h000;
    rom[9641 ] = 12'h000;
    rom[9642 ] = 12'h000;
    rom[9643 ] = 12'h000;
    rom[9644 ] = 12'h000;
    rom[9645 ] = 12'h000;
    rom[9646 ] = 12'h000;
    rom[9647 ] = 12'h000;
    rom[9648 ] = 12'h000;
    rom[9649 ] = 12'h000;
    rom[9650 ] = 12'h000;
    rom[9651 ] = 12'h000;
    rom[9652 ] = 12'h000;
    rom[9653 ] = 12'h000;
    rom[9654 ] = 12'h000;
    rom[9655 ] = 12'h000;
    rom[9656 ] = 12'h3a2;
    rom[9657 ] = 12'h3a2;
    rom[9658 ] = 12'h3a2;
    rom[9659 ] = 12'h3a2;
    rom[9660 ] = 12'h3a2;
    rom[9661 ] = 12'h3a2;
    rom[9662 ] = 12'h3a2;
    rom[9663 ] = 12'h3a2;
    rom[9664 ] = 12'h3a2;
    rom[9665 ] = 12'h3a2;
    rom[9666 ] = 12'h3a2;
    rom[9667 ] = 12'h3a2;
    rom[9668 ] = 12'h3a2;
    rom[9669 ] = 12'h3a2;
    rom[9670 ] = 12'h3a2;
    rom[9671 ] = 12'h000;
    rom[9672 ] = 12'h000;
    rom[9673 ] = 12'h000;
    rom[9674 ] = 12'h000;
    rom[9675 ] = 12'h000;
    rom[9676 ] = 12'h000;
    rom[9677 ] = 12'h000;
    rom[9678 ] = 12'h000;
    rom[9679 ] = 12'h000;
    rom[9680 ] = 12'h000;
    rom[9681 ] = 12'h000;
    rom[9682 ] = 12'h000;
    rom[9683 ] = 12'h000;
    rom[9684 ] = 12'h000;
    rom[9685 ] = 12'h000;
    rom[9686 ] = 12'h000;
    rom[9687 ] = 12'h000;
    rom[9688 ] = 12'h000;
    rom[9689 ] = 12'h000;
    rom[9690 ] = 12'h000;
    rom[9691 ] = 12'h000;
    rom[9692 ] = 12'h000;
    rom[9693 ] = 12'h000;
    rom[9694 ] = 12'h000;
    rom[9695 ] = 12'h000;
    rom[9696 ] = 12'h000;
    rom[9697 ] = 12'h000;
    rom[9698 ] = 12'h000;
    rom[9699 ] = 12'h000;
    rom[9700 ] = 12'h000;
    rom[9701 ] = 12'h000;
    rom[9702 ] = 12'h000;
    rom[9703 ] = 12'h000;
    rom[9704 ] = 12'h000;
    rom[9705 ] = 12'h000;
    rom[9706 ] = 12'h000;
    rom[9707 ] = 12'h000;
    rom[9708 ] = 12'h000;
    rom[9709 ] = 12'h000;
    rom[9710 ] = 12'h000;
    rom[9711 ] = 12'h000;
    rom[9712 ] = 12'h3a2;
    rom[9713 ] = 12'h3a2;
    rom[9714 ] = 12'h3a2;
    rom[9715 ] = 12'h3a2;
    rom[9716 ] = 12'h3a2;
    rom[9717 ] = 12'h3a2;
    rom[9718 ] = 12'h3a2;
    rom[9719 ] = 12'h3a2;
    rom[9720 ] = 12'h3a2;
    rom[9721 ] = 12'h3a2;
    rom[9722 ] = 12'h3a2;
    rom[9723 ] = 12'h3a2;
    rom[9724 ] = 12'h3a2;
    rom[9725 ] = 12'h3a2;
    rom[9726 ] = 12'h3a2;
    rom[9727 ] = 12'h000;
    rom[9728 ] = 12'h000;
    rom[9729 ] = 12'h3db;
    rom[9730 ] = 12'h3db;
    rom[9731 ] = 12'h2db;
    rom[9732 ] = 12'h2db;
    rom[9733 ] = 12'h2db;
    rom[9734 ] = 12'h2db;
    rom[9735 ] = 12'h2db;
    rom[9736 ] = 12'h2db;
    rom[9737 ] = 12'h2db;
    rom[9738 ] = 12'h2db;
    rom[9739 ] = 12'h2db;
    rom[9740 ] = 12'h2db;
    rom[9741 ] = 12'h2dc;
    rom[9742 ] = 12'h2dc;
    rom[9743 ] = 12'h2dc;
    rom[9744 ] = 12'h000;
    rom[9745 ] = 12'h000;
    rom[9746 ] = 12'h000;
    rom[9747 ] = 12'h000;
    rom[9748 ] = 12'h000;
    rom[9749 ] = 12'h000;
    rom[9750 ] = 12'h000;
    rom[9751 ] = 12'h000;
    rom[9752 ] = 12'h000;
    rom[9753 ] = 12'h000;
    rom[9754 ] = 12'h000;
    rom[9755 ] = 12'h000;
    rom[9756 ] = 12'h000;
    rom[9757 ] = 12'h000;
    rom[9758 ] = 12'h000;
    rom[9759 ] = 12'h000;
    rom[9760 ] = 12'h000;
    rom[9761 ] = 12'h000;
    rom[9762 ] = 12'h000;
    rom[9763 ] = 12'h000;
    rom[9764 ] = 12'h000;
    rom[9765 ] = 12'h000;
    rom[9766 ] = 12'h000;
    rom[9767 ] = 12'h000;
    rom[9768 ] = 12'h000;
    rom[9769 ] = 12'h000;
    rom[9770 ] = 12'h000;
    rom[9771 ] = 12'h000;
    rom[9772 ] = 12'h000;
    rom[9773 ] = 12'h000;
    rom[9774 ] = 12'h000;
    rom[9775 ] = 12'h000;
    rom[9776 ] = 12'h000;
    rom[9777 ] = 12'h000;
    rom[9778 ] = 12'h000;
    rom[9779 ] = 12'h000;
    rom[9780 ] = 12'h000;
    rom[9781 ] = 12'h000;
    rom[9782 ] = 12'h000;
    rom[9783 ] = 12'h000;
    rom[9784 ] = 12'h000;
    rom[9785 ] = 12'h3a2;
    rom[9786 ] = 12'h3a2;
    rom[9787 ] = 12'h3a2;
    rom[9788 ] = 12'h3a2;
    rom[9789 ] = 12'h3a2;
    rom[9790 ] = 12'h3a2;
    rom[9791 ] = 12'h3a2;
    rom[9792 ] = 12'h3a2;
    rom[9793 ] = 12'h3a2;
    rom[9794 ] = 12'h3a2;
    rom[9795 ] = 12'h3a2;
    rom[9796 ] = 12'h3a2;
    rom[9797 ] = 12'h3a2;
    rom[9798 ] = 12'h000;
    rom[9799 ] = 12'h000;
    rom[9800 ] = 12'h000;
    rom[9801 ] = 12'h000;
    rom[9802 ] = 12'h000;
    rom[9803 ] = 12'h000;
    rom[9804 ] = 12'h000;
    rom[9805 ] = 12'h000;
    rom[9806 ] = 12'h000;
    rom[9807 ] = 12'h000;
    rom[9808 ] = 12'h000;
    rom[9809 ] = 12'h000;
    rom[9810 ] = 12'h000;
    rom[9811 ] = 12'h000;
    rom[9812 ] = 12'h000;
    rom[9813 ] = 12'h000;
    rom[9814 ] = 12'h000;
    rom[9815 ] = 12'h000;
    rom[9816 ] = 12'h000;
    rom[9817 ] = 12'h000;
    rom[9818 ] = 12'h000;
    rom[9819 ] = 12'h000;
    rom[9820 ] = 12'h000;
    rom[9821 ] = 12'h000;
    rom[9822 ] = 12'h000;
    rom[9823 ] = 12'h000;
    rom[9824 ] = 12'h000;
    rom[9825 ] = 12'h000;
    rom[9826 ] = 12'h000;
    rom[9827 ] = 12'h000;
    rom[9828 ] = 12'h000;
    rom[9829 ] = 12'h000;
    rom[9830 ] = 12'h000;
    rom[9831 ] = 12'h000;
    rom[9832 ] = 12'h000;
    rom[9833 ] = 12'h000;
    rom[9834 ] = 12'h000;
    rom[9835 ] = 12'h000;
    rom[9836 ] = 12'h000;
    rom[9837 ] = 12'h000;
    rom[9838 ] = 12'h000;
    rom[9839 ] = 12'h000;
    rom[9840 ] = 12'h3a2;
    rom[9841 ] = 12'h3a2;
    rom[9842 ] = 12'h3a2;
    rom[9843 ] = 12'h3a2;
    rom[9844 ] = 12'h3a2;
    rom[9845 ] = 12'h3a2;
    rom[9846 ] = 12'h3a2;
    rom[9847 ] = 12'h3a2;
    rom[9848 ] = 12'h3a2;
    rom[9849 ] = 12'h3a2;
    rom[9850 ] = 12'h3a2;
    rom[9851 ] = 12'h3a2;
    rom[9852 ] = 12'h3a2;
    rom[9853 ] = 12'h3a2;
    rom[9854 ] = 12'h3a2;
    rom[9855 ] = 12'h000;
    rom[9856 ] = 12'h000;
    rom[9857 ] = 12'h2db;
    rom[9858 ] = 12'h2db;
    rom[9859 ] = 12'h2db;
    rom[9860 ] = 12'h2db;
    rom[9861 ] = 12'h2db;
    rom[9862 ] = 12'h2db;
    rom[9863 ] = 12'h2db;
    rom[9864 ] = 12'h2db;
    rom[9865 ] = 12'h2db;
    rom[9866 ] = 12'h2dc;
    rom[9867 ] = 12'h2dc;
    rom[9868 ] = 12'h2dc;
    rom[9869 ] = 12'h2dc;
    rom[9870 ] = 12'h2dc;
    rom[9871 ] = 12'h2dc;
    rom[9872 ] = 12'h2dc;
    rom[9873 ] = 12'h000;
    rom[9874 ] = 12'h000;
    rom[9875 ] = 12'h000;
    rom[9876 ] = 12'h000;
    rom[9877 ] = 12'h000;
    rom[9878 ] = 12'h000;
    rom[9879 ] = 12'h000;
    rom[9880 ] = 12'h000;
    rom[9881 ] = 12'h000;
    rom[9882 ] = 12'h000;
    rom[9883 ] = 12'h000;
    rom[9884 ] = 12'h000;
    rom[9885 ] = 12'h000;
    rom[9886 ] = 12'h000;
    rom[9887 ] = 12'h000;
    rom[9888 ] = 12'h000;
    rom[9889 ] = 12'h000;
    rom[9890 ] = 12'h000;
    rom[9891 ] = 12'h000;
    rom[9892 ] = 12'h000;
    rom[9893 ] = 12'h000;
    rom[9894 ] = 12'h000;
    rom[9895 ] = 12'h000;
    rom[9896 ] = 12'h000;
    rom[9897 ] = 12'h000;
    rom[9898 ] = 12'h000;
    rom[9899 ] = 12'h000;
    rom[9900 ] = 12'h000;
    rom[9901 ] = 12'h000;
    rom[9902 ] = 12'h000;
    rom[9903 ] = 12'h000;
    rom[9904 ] = 12'h000;
    rom[9905 ] = 12'h000;
    rom[9906 ] = 12'h000;
    rom[9907 ] = 12'h000;
    rom[9908 ] = 12'h000;
    rom[9909 ] = 12'h000;
    rom[9910 ] = 12'h000;
    rom[9911 ] = 12'h000;
    rom[9912 ] = 12'h000;
    rom[9913 ] = 12'h000;
    rom[9914 ] = 12'h000;
    rom[9915 ] = 12'h3a2;
    rom[9916 ] = 12'h3a2;
    rom[9917 ] = 12'h3a2;
    rom[9918 ] = 12'h3a2;
    rom[9919 ] = 12'h3a2;
    rom[9920 ] = 12'h3a2;
    rom[9921 ] = 12'h3a2;
    rom[9922 ] = 12'h3a2;
    rom[9923 ] = 12'h3a2;
    rom[9924 ] = 12'h3a2;
    rom[9925 ] = 12'h000;
    rom[9926 ] = 12'h000;
    rom[9927 ] = 12'h000;
    rom[9928 ] = 12'h000;
    rom[9929 ] = 12'h000;
    rom[9930 ] = 12'h000;
    rom[9931 ] = 12'h000;
    rom[9932 ] = 12'h000;
    rom[9933 ] = 12'h000;
    rom[9934 ] = 12'h000;
    rom[9935 ] = 12'h000;
    rom[9936 ] = 12'h000;
    rom[9937 ] = 12'h000;
    rom[9938 ] = 12'h000;
    rom[9939 ] = 12'h000;
    rom[9940 ] = 12'h000;
    rom[9941 ] = 12'h000;
    rom[9942 ] = 12'h000;
    rom[9943 ] = 12'h000;
    rom[9944 ] = 12'h000;
    rom[9945 ] = 12'h000;
    rom[9946 ] = 12'h000;
    rom[9947 ] = 12'h000;
    rom[9948 ] = 12'h000;
    rom[9949 ] = 12'h000;
    rom[9950 ] = 12'h000;
    rom[9951 ] = 12'h000;
    rom[9952 ] = 12'h000;
    rom[9953 ] = 12'h000;
    rom[9954 ] = 12'h000;
    rom[9955 ] = 12'h000;
    rom[9956 ] = 12'h000;
    rom[9957 ] = 12'h000;
    rom[9958 ] = 12'h000;
    rom[9959 ] = 12'h000;
    rom[9960 ] = 12'h000;
    rom[9961 ] = 12'h000;
    rom[9962 ] = 12'h000;
    rom[9963 ] = 12'h000;
    rom[9964 ] = 12'h000;
    rom[9965 ] = 12'h000;
    rom[9966 ] = 12'h000;
    rom[9967 ] = 12'h3a2;
    rom[9968 ] = 12'h3a2;
    rom[9969 ] = 12'h3a2;
    rom[9970 ] = 12'h3a2;
    rom[9971 ] = 12'h3a2;
    rom[9972 ] = 12'h3a2;
    rom[9973 ] = 12'h3a2;
    rom[9974 ] = 12'h3a2;
    rom[9975 ] = 12'h3a2;
    rom[9976 ] = 12'h3a2;
    rom[9977 ] = 12'h3a2;
    rom[9978 ] = 12'h3a2;
    rom[9979 ] = 12'h3a2;
    rom[9980 ] = 12'h3a2;
    rom[9981 ] = 12'h3a2;
    rom[9982 ] = 12'h3a2;
    rom[9983 ] = 12'h000;
    rom[9984 ] = 12'h000;
    rom[9985 ] = 12'h000;
    rom[9986 ] = 12'h2db;
    rom[9987 ] = 12'h2db;
    rom[9988 ] = 12'h2db;
    rom[9989 ] = 12'h2db;
    rom[9990 ] = 12'h2db;
    rom[9991 ] = 12'h2dc;
    rom[9992 ] = 12'h2dc;
    rom[9993 ] = 12'h2dc;
    rom[9994 ] = 12'h2dc;
    rom[9995 ] = 12'h2dc;
    rom[9996 ] = 12'h2dc;
    rom[9997 ] = 12'h2dc;
    rom[9998 ] = 12'h2dc;
    rom[9999 ] = 12'h2dc;
    rom[10000] = 12'h2dc;
    rom[10001] = 12'h000;
    rom[10002] = 12'h000;
    rom[10003] = 12'h000;
    rom[10004] = 12'h000;
    rom[10005] = 12'h000;
    rom[10006] = 12'h000;
    rom[10007] = 12'h000;
    rom[10008] = 12'h000;
    rom[10009] = 12'h000;
    rom[10010] = 12'h000;
    rom[10011] = 12'h000;
    rom[10012] = 12'h000;
    rom[10013] = 12'h000;
    rom[10014] = 12'h000;
    rom[10015] = 12'h000;
    rom[10016] = 12'h000;
    rom[10017] = 12'h000;
    rom[10018] = 12'h000;
    rom[10019] = 12'h000;
    rom[10020] = 12'h000;
    rom[10021] = 12'h000;
    rom[10022] = 12'h000;
    rom[10023] = 12'h000;
    rom[10024] = 12'h000;
    rom[10025] = 12'h000;
    rom[10026] = 12'h000;
    rom[10027] = 12'h000;
    rom[10028] = 12'h000;
    rom[10029] = 12'h000;
    rom[10030] = 12'h000;
    rom[10031] = 12'h000;
    rom[10032] = 12'h000;
    rom[10033] = 12'h000;
    rom[10034] = 12'h000;
    rom[10035] = 12'h000;
    rom[10036] = 12'h000;
    rom[10037] = 12'h000;
    rom[10038] = 12'h000;
    rom[10039] = 12'h000;
    rom[10040] = 12'h000;
    rom[10041] = 12'h000;
    rom[10042] = 12'h000;
    rom[10043] = 12'h000;
    rom[10044] = 12'h3a2;
    rom[10045] = 12'h3a2;
    rom[10046] = 12'h3a2;
    rom[10047] = 12'h3a2;
    rom[10048] = 12'h3a2;
    rom[10049] = 12'h3a2;
    rom[10050] = 12'h3a2;
    rom[10051] = 12'h000;
    rom[10052] = 12'h000;
    rom[10053] = 12'h000;
    rom[10054] = 12'h000;
    rom[10055] = 12'h000;
    rom[10056] = 12'h000;
    rom[10057] = 12'h000;
    rom[10058] = 12'h000;
    rom[10059] = 12'h000;
    rom[10060] = 12'h000;
    rom[10061] = 12'h000;
    rom[10062] = 12'h000;
    rom[10063] = 12'h000;
    rom[10064] = 12'h000;
    rom[10065] = 12'h000;
    rom[10066] = 12'h000;
    rom[10067] = 12'h000;
    rom[10068] = 12'h000;
    rom[10069] = 12'h000;
    rom[10070] = 12'h000;
    rom[10071] = 12'h000;
    rom[10072] = 12'h000;
    rom[10073] = 12'h000;
    rom[10074] = 12'h000;
    rom[10075] = 12'h000;
    rom[10076] = 12'h000;
    rom[10077] = 12'h000;
    rom[10078] = 12'h000;
    rom[10079] = 12'h000;
    rom[10080] = 12'h000;
    rom[10081] = 12'h000;
    rom[10082] = 12'h000;
    rom[10083] = 12'h000;
    rom[10084] = 12'h000;
    rom[10085] = 12'h000;
    rom[10086] = 12'h000;
    rom[10087] = 12'h000;
    rom[10088] = 12'h000;
    rom[10089] = 12'h000;
    rom[10090] = 12'h000;
    rom[10091] = 12'h000;
    rom[10092] = 12'h000;
    rom[10093] = 12'h000;
    rom[10094] = 12'h000;
    rom[10095] = 12'h3a2;
    rom[10096] = 12'h3a2;
    rom[10097] = 12'h3a2;
    rom[10098] = 12'h3a2;
    rom[10099] = 12'h3a2;
    rom[10100] = 12'h3a2;
    rom[10101] = 12'h3a2;
    rom[10102] = 12'h3a2;
    rom[10103] = 12'h3a2;
    rom[10104] = 12'h3a2;
    rom[10105] = 12'h3a2;
    rom[10106] = 12'h3a2;
    rom[10107] = 12'h3a2;
    rom[10108] = 12'h3a2;
    rom[10109] = 12'h3a2;
    rom[10110] = 12'h000;
    rom[10111] = 12'h000;
    rom[10112] = 12'h000;
    rom[10113] = 12'h000;
    rom[10114] = 12'h2db;
    rom[10115] = 12'h2db;
    rom[10116] = 12'h2dc;
    rom[10117] = 12'h2dc;
    rom[10118] = 12'h2dc;
    rom[10119] = 12'h2dc;
    rom[10120] = 12'h2dc;
    rom[10121] = 12'h2dc;
    rom[10122] = 12'h2dc;
    rom[10123] = 12'h2dc;
    rom[10124] = 12'h2dc;
    rom[10125] = 12'h2dc;
    rom[10126] = 12'h2dc;
    rom[10127] = 12'h2dc;
    rom[10128] = 12'h2dc;
    rom[10129] = 12'h000;
    rom[10130] = 12'h000;
    rom[10131] = 12'h000;
    rom[10132] = 12'h000;
    rom[10133] = 12'h000;
    rom[10134] = 12'h000;
    rom[10135] = 12'h000;
    rom[10136] = 12'h000;
    rom[10137] = 12'h000;
    rom[10138] = 12'h000;
    rom[10139] = 12'h000;
    rom[10140] = 12'h000;
    rom[10141] = 12'h000;
    rom[10142] = 12'h000;
    rom[10143] = 12'h000;
    rom[10144] = 12'h000;
    rom[10145] = 12'h000;
    rom[10146] = 12'h000;
    rom[10147] = 12'h000;
    rom[10148] = 12'h000;
    rom[10149] = 12'h000;
    rom[10150] = 12'h000;
    rom[10151] = 12'h000;
    rom[10152] = 12'h000;
    rom[10153] = 12'h000;
    rom[10154] = 12'h000;
    rom[10155] = 12'h000;
    rom[10156] = 12'h000;
    rom[10157] = 12'h000;
    rom[10158] = 12'h000;
    rom[10159] = 12'h000;
    rom[10160] = 12'h000;
    rom[10161] = 12'h000;
    rom[10162] = 12'h000;
    rom[10163] = 12'h000;
    rom[10164] = 12'h000;
    rom[10165] = 12'h000;
    rom[10166] = 12'h000;
    rom[10167] = 12'h000;
    rom[10168] = 12'h000;
    rom[10169] = 12'h000;
    rom[10170] = 12'h000;
    rom[10171] = 12'h000;
    rom[10172] = 12'h000;
    rom[10173] = 12'h000;
    rom[10174] = 12'h3a2;
    rom[10175] = 12'h3a2;
    rom[10176] = 12'h3a2;
    rom[10177] = 12'h3a2;
    rom[10178] = 12'h000;
    rom[10179] = 12'h000;
    rom[10180] = 12'h000;
    rom[10181] = 12'h000;
    rom[10182] = 12'h000;
    rom[10183] = 12'h000;
    rom[10184] = 12'h000;
    rom[10185] = 12'h000;
    rom[10186] = 12'h000;
    rom[10187] = 12'h000;
    rom[10188] = 12'h000;
    rom[10189] = 12'h000;
    rom[10190] = 12'h000;
    rom[10191] = 12'h000;
    rom[10192] = 12'h000;
    rom[10193] = 12'h000;
    rom[10194] = 12'h000;
    rom[10195] = 12'h000;
    rom[10196] = 12'h000;
    rom[10197] = 12'h000;
    rom[10198] = 12'h000;
    rom[10199] = 12'h000;
    rom[10200] = 12'h000;
    rom[10201] = 12'h000;
    rom[10202] = 12'h000;
    rom[10203] = 12'h000;
    rom[10204] = 12'h000;
    rom[10205] = 12'h000;
    rom[10206] = 12'h000;
    rom[10207] = 12'h000;
    rom[10208] = 12'h000;
    rom[10209] = 12'h000;
    rom[10210] = 12'h000;
    rom[10211] = 12'h000;
    rom[10212] = 12'h000;
    rom[10213] = 12'h000;
    rom[10214] = 12'h000;
    rom[10215] = 12'h000;
    rom[10216] = 12'h000;
    rom[10217] = 12'h000;
    rom[10218] = 12'h000;
    rom[10219] = 12'h000;
    rom[10220] = 12'h000;
    rom[10221] = 12'h000;
    rom[10222] = 12'h000;
    rom[10223] = 12'h3a2;
    rom[10224] = 12'h3a2;
    rom[10225] = 12'h3a2;
    rom[10226] = 12'h3a2;
    rom[10227] = 12'h3a2;
    rom[10228] = 12'h3a2;
    rom[10229] = 12'h3a2;
    rom[10230] = 12'h3a2;
    rom[10231] = 12'h3a2;
    rom[10232] = 12'h3a2;
    rom[10233] = 12'h3a2;
    rom[10234] = 12'h3a2;
    rom[10235] = 12'h3a2;
    rom[10236] = 12'h3a2;
    rom[10237] = 12'h3a2;
    rom[10238] = 12'h000;
    rom[10239] = 12'h000;
    rom[10240] = 12'h000;
    rom[10241] = 12'h000;
    rom[10242] = 12'h2dc;
    rom[10243] = 12'h2dc;
    rom[10244] = 12'h2dc;
    rom[10245] = 12'h2dc;
    rom[10246] = 12'h2dc;
    rom[10247] = 12'h2dc;
    rom[10248] = 12'h2dc;
    rom[10249] = 12'h2dc;
    rom[10250] = 12'h2dc;
    rom[10251] = 12'h2dc;
    rom[10252] = 12'h2dc;
    rom[10253] = 12'h2dc;
    rom[10254] = 12'h2dc;
    rom[10255] = 12'h2dc;
    rom[10256] = 12'h2dc;
    rom[10257] = 12'h2dc;
    rom[10258] = 12'h000;
    rom[10259] = 12'h000;
    rom[10260] = 12'h000;
    rom[10261] = 12'h000;
    rom[10262] = 12'h000;
    rom[10263] = 12'h000;
    rom[10264] = 12'h000;
    rom[10265] = 12'h000;
    rom[10266] = 12'h000;
    rom[10267] = 12'h000;
    rom[10268] = 12'h000;
    rom[10269] = 12'h000;
    rom[10270] = 12'h000;
    rom[10271] = 12'h000;
    rom[10272] = 12'h000;
    rom[10273] = 12'h000;
    rom[10274] = 12'h000;
    rom[10275] = 12'h000;
    rom[10276] = 12'h000;
    rom[10277] = 12'h000;
    rom[10278] = 12'h000;
    rom[10279] = 12'h000;
    rom[10280] = 12'h000;
    rom[10281] = 12'h000;
    rom[10282] = 12'h000;
    rom[10283] = 12'h000;
    rom[10284] = 12'h000;
    rom[10285] = 12'h000;
    rom[10286] = 12'h000;
    rom[10287] = 12'h000;
    rom[10288] = 12'h000;
    rom[10289] = 12'h000;
    rom[10290] = 12'h000;
    rom[10291] = 12'h000;
    rom[10292] = 12'h000;
    rom[10293] = 12'h000;
    rom[10294] = 12'h000;
    rom[10295] = 12'h000;
    rom[10296] = 12'h000;
    rom[10297] = 12'h000;
    rom[10298] = 12'h000;
    rom[10299] = 12'h000;
    rom[10300] = 12'h000;
    rom[10301] = 12'h000;
    rom[10302] = 12'h000;
    rom[10303] = 12'h000;
    rom[10304] = 12'h393;
    rom[10305] = 12'h000;
    rom[10306] = 12'h000;
    rom[10307] = 12'h000;
    rom[10308] = 12'h000;
    rom[10309] = 12'h000;
    rom[10310] = 12'h000;
    rom[10311] = 12'h000;
    rom[10312] = 12'h000;
    rom[10313] = 12'h000;
    rom[10314] = 12'h000;
    rom[10315] = 12'h000;
    rom[10316] = 12'h000;
    rom[10317] = 12'h000;
    rom[10318] = 12'h000;
    rom[10319] = 12'h000;
    rom[10320] = 12'h000;
    rom[10321] = 12'h000;
    rom[10322] = 12'h000;
    rom[10323] = 12'h000;
    rom[10324] = 12'h000;
    rom[10325] = 12'h000;
    rom[10326] = 12'h000;
    rom[10327] = 12'h000;
    rom[10328] = 12'h000;
    rom[10329] = 12'h000;
    rom[10330] = 12'h000;
    rom[10331] = 12'h000;
    rom[10332] = 12'h000;
    rom[10333] = 12'h000;
    rom[10334] = 12'h000;
    rom[10335] = 12'h000;
    rom[10336] = 12'h000;
    rom[10337] = 12'h000;
    rom[10338] = 12'h000;
    rom[10339] = 12'h000;
    rom[10340] = 12'h000;
    rom[10341] = 12'h000;
    rom[10342] = 12'h000;
    rom[10343] = 12'h000;
    rom[10344] = 12'h000;
    rom[10345] = 12'h000;
    rom[10346] = 12'h000;
    rom[10347] = 12'h000;
    rom[10348] = 12'h000;
    rom[10349] = 12'h000;
    rom[10350] = 12'h3a2;
    rom[10351] = 12'h3a2;
    rom[10352] = 12'h3a2;
    rom[10353] = 12'h3a2;
    rom[10354] = 12'h3a2;
    rom[10355] = 12'h3a2;
    rom[10356] = 12'h3a2;
    rom[10357] = 12'h3a2;
    rom[10358] = 12'h3a2;
    rom[10359] = 12'h3a2;
    rom[10360] = 12'h3a2;
    rom[10361] = 12'h3a2;
    rom[10362] = 12'h3a2;
    rom[10363] = 12'h3a2;
    rom[10364] = 12'h3a2;
    rom[10365] = 12'h3a2;
    rom[10366] = 12'h000;
    rom[10367] = 12'h000;
    rom[10368] = 12'h000;
    rom[10369] = 12'h000;
    rom[10370] = 12'h2dc;
    rom[10371] = 12'h2dc;
    rom[10372] = 12'h2dc;
    rom[10373] = 12'h2dc;
    rom[10374] = 12'h2dc;
    rom[10375] = 12'h2dc;
    rom[10376] = 12'h2dc;
    rom[10377] = 12'h2dc;
    rom[10378] = 12'h2dc;
    rom[10379] = 12'h2dc;
    rom[10380] = 12'h2dc;
    rom[10381] = 12'h2dc;
    rom[10382] = 12'h2dc;
    rom[10383] = 12'h2dc;
    rom[10384] = 12'h2dc;
    rom[10385] = 12'h2dc;
    rom[10386] = 12'h000;
    rom[10387] = 12'h000;
    rom[10388] = 12'h000;
    rom[10389] = 12'h000;
    rom[10390] = 12'h000;
    rom[10391] = 12'h000;
    rom[10392] = 12'h000;
    rom[10393] = 12'h000;
    rom[10394] = 12'h000;
    rom[10395] = 12'h000;
    rom[10396] = 12'h000;
    rom[10397] = 12'h000;
    rom[10398] = 12'h000;
    rom[10399] = 12'h000;
    rom[10400] = 12'h000;
    rom[10401] = 12'h000;
    rom[10402] = 12'h000;
    rom[10403] = 12'h000;
    rom[10404] = 12'h000;
    rom[10405] = 12'h000;
    rom[10406] = 12'h000;
    rom[10407] = 12'h000;
    rom[10408] = 12'h000;
    rom[10409] = 12'h000;
    rom[10410] = 12'h000;
    rom[10411] = 12'h000;
    rom[10412] = 12'h000;
    rom[10413] = 12'h000;
    rom[10414] = 12'h000;
    rom[10415] = 12'h000;
    rom[10416] = 12'h000;
    rom[10417] = 12'h000;
    rom[10418] = 12'h000;
    rom[10419] = 12'h000;
    rom[10420] = 12'h000;
    rom[10421] = 12'h000;
    rom[10422] = 12'h000;
    rom[10423] = 12'h000;
    rom[10424] = 12'h000;
    rom[10425] = 12'h000;
    rom[10426] = 12'h000;
    rom[10427] = 12'h000;
    rom[10428] = 12'h000;
    rom[10429] = 12'h000;
    rom[10430] = 12'h000;
    rom[10431] = 12'h000;
    rom[10432] = 12'h000;
    rom[10433] = 12'h000;
    rom[10434] = 12'h000;
    rom[10435] = 12'h000;
    rom[10436] = 12'h000;
    rom[10437] = 12'h000;
    rom[10438] = 12'h000;
    rom[10439] = 12'h000;
    rom[10440] = 12'h000;
    rom[10441] = 12'h000;
    rom[10442] = 12'h000;
    rom[10443] = 12'h000;
    rom[10444] = 12'h000;
    rom[10445] = 12'h000;
    rom[10446] = 12'h000;
    rom[10447] = 12'h000;
    rom[10448] = 12'h000;
    rom[10449] = 12'h000;
    rom[10450] = 12'h000;
    rom[10451] = 12'h000;
    rom[10452] = 12'h000;
    rom[10453] = 12'h000;
    rom[10454] = 12'h000;
    rom[10455] = 12'h000;
    rom[10456] = 12'h000;
    rom[10457] = 12'h000;
    rom[10458] = 12'h000;
    rom[10459] = 12'h000;
    rom[10460] = 12'h000;
    rom[10461] = 12'h000;
    rom[10462] = 12'h000;
    rom[10463] = 12'h000;
    rom[10464] = 12'h000;
    rom[10465] = 12'h000;
    rom[10466] = 12'h000;
    rom[10467] = 12'h000;
    rom[10468] = 12'h000;
    rom[10469] = 12'h000;
    rom[10470] = 12'h000;
    rom[10471] = 12'h000;
    rom[10472] = 12'h000;
    rom[10473] = 12'h000;
    rom[10474] = 12'h000;
    rom[10475] = 12'h000;
    rom[10476] = 12'h000;
    rom[10477] = 12'h000;
    rom[10478] = 12'h3a2;
    rom[10479] = 12'h3a2;
    rom[10480] = 12'h3a2;
    rom[10481] = 12'h3a2;
    rom[10482] = 12'h3a2;
    rom[10483] = 12'h3a2;
    rom[10484] = 12'h3a2;
    rom[10485] = 12'h3a2;
    rom[10486] = 12'h3a2;
    rom[10487] = 12'h3a2;
    rom[10488] = 12'h3a2;
    rom[10489] = 12'h3a2;
    rom[10490] = 12'h3a2;
    rom[10491] = 12'h3a2;
    rom[10492] = 12'h3a2;
    rom[10493] = 12'h392;
    rom[10494] = 12'h000;
    rom[10495] = 12'h000;
    rom[10496] = 12'h000;
    rom[10497] = 12'h000;
    rom[10498] = 12'h000;
    rom[10499] = 12'h2dc;
    rom[10500] = 12'h2dc;
    rom[10501] = 12'h2dc;
    rom[10502] = 12'h2dc;
    rom[10503] = 12'h2dc;
    rom[10504] = 12'h2dc;
    rom[10505] = 12'h2dc;
    rom[10506] = 12'h2dc;
    rom[10507] = 12'h2dc;
    rom[10508] = 12'h2dc;
    rom[10509] = 12'h2dc;
    rom[10510] = 12'h2dc;
    rom[10511] = 12'h2dd;
    rom[10512] = 12'h2dd;
    rom[10513] = 12'h2dd;
    rom[10514] = 12'h3cc;
    rom[10515] = 12'h000;
    rom[10516] = 12'h000;
    rom[10517] = 12'h000;
    rom[10518] = 12'h000;
    rom[10519] = 12'h000;
    rom[10520] = 12'h000;
    rom[10521] = 12'h000;
    rom[10522] = 12'h000;
    rom[10523] = 12'h000;
    rom[10524] = 12'h000;
    rom[10525] = 12'h000;
    rom[10526] = 12'h000;
    rom[10527] = 12'h000;
    rom[10528] = 12'h000;
    rom[10529] = 12'h000;
    rom[10530] = 12'h000;
    rom[10531] = 12'h000;
    rom[10532] = 12'h000;
    rom[10533] = 12'h000;
    rom[10534] = 12'h000;
    rom[10535] = 12'h000;
    rom[10536] = 12'h000;
    rom[10537] = 12'h000;
    rom[10538] = 12'h000;
    rom[10539] = 12'h000;
    rom[10540] = 12'h000;
    rom[10541] = 12'h000;
    rom[10542] = 12'h000;
    rom[10543] = 12'h000;
    rom[10544] = 12'h000;
    rom[10545] = 12'h000;
    rom[10546] = 12'h000;
    rom[10547] = 12'h000;
    rom[10548] = 12'h000;
    rom[10549] = 12'h000;
    rom[10550] = 12'h000;
    rom[10551] = 12'h000;
    rom[10552] = 12'h000;
    rom[10553] = 12'h000;
    rom[10554] = 12'h000;
    rom[10555] = 12'h000;
    rom[10556] = 12'h000;
    rom[10557] = 12'h000;
    rom[10558] = 12'h000;
    rom[10559] = 12'h000;
    rom[10560] = 12'h000;
    rom[10561] = 12'h000;
    rom[10562] = 12'h000;
    rom[10563] = 12'h000;
    rom[10564] = 12'h000;
    rom[10565] = 12'h000;
    rom[10566] = 12'h000;
    rom[10567] = 12'h000;
    rom[10568] = 12'h000;
    rom[10569] = 12'h000;
    rom[10570] = 12'h000;
    rom[10571] = 12'h000;
    rom[10572] = 12'h000;
    rom[10573] = 12'h000;
    rom[10574] = 12'h000;
    rom[10575] = 12'h000;
    rom[10576] = 12'h000;
    rom[10577] = 12'h000;
    rom[10578] = 12'h000;
    rom[10579] = 12'h000;
    rom[10580] = 12'h000;
    rom[10581] = 12'h000;
    rom[10582] = 12'h000;
    rom[10583] = 12'h000;
    rom[10584] = 12'h000;
    rom[10585] = 12'h000;
    rom[10586] = 12'h000;
    rom[10587] = 12'h000;
    rom[10588] = 12'h000;
    rom[10589] = 12'h000;
    rom[10590] = 12'h000;
    rom[10591] = 12'h000;
    rom[10592] = 12'h000;
    rom[10593] = 12'h000;
    rom[10594] = 12'h000;
    rom[10595] = 12'h000;
    rom[10596] = 12'h000;
    rom[10597] = 12'h000;
    rom[10598] = 12'h000;
    rom[10599] = 12'h000;
    rom[10600] = 12'h000;
    rom[10601] = 12'h000;
    rom[10602] = 12'h000;
    rom[10603] = 12'h000;
    rom[10604] = 12'h000;
    rom[10605] = 12'h492;
    rom[10606] = 12'h3a2;
    rom[10607] = 12'h3a2;
    rom[10608] = 12'h3a2;
    rom[10609] = 12'h3a2;
    rom[10610] = 12'h3a2;
    rom[10611] = 12'h3a2;
    rom[10612] = 12'h3a2;
    rom[10613] = 12'h3a2;
    rom[10614] = 12'h3a2;
    rom[10615] = 12'h3a2;
    rom[10616] = 12'h3a2;
    rom[10617] = 12'h3a2;
    rom[10618] = 12'h3a2;
    rom[10619] = 12'h3a2;
    rom[10620] = 12'h3a2;
    rom[10621] = 12'h000;
    rom[10622] = 12'h000;
    rom[10623] = 12'h000;
    rom[10624] = 12'h000;
    rom[10625] = 12'h000;
    rom[10626] = 12'h000;
    rom[10627] = 12'h2dc;
    rom[10628] = 12'h2dc;
    rom[10629] = 12'h2dc;
    rom[10630] = 12'h2dc;
    rom[10631] = 12'h2dc;
    rom[10632] = 12'h2dc;
    rom[10633] = 12'h2dc;
    rom[10634] = 12'h2dc;
    rom[10635] = 12'h2dc;
    rom[10636] = 12'h2dd;
    rom[10637] = 12'h2dd;
    rom[10638] = 12'h2dd;
    rom[10639] = 12'h2dd;
    rom[10640] = 12'h2dd;
    rom[10641] = 12'h2dd;
    rom[10642] = 12'h2dd;
    rom[10643] = 12'h000;
    rom[10644] = 12'h000;
    rom[10645] = 12'h000;
    rom[10646] = 12'h000;
    rom[10647] = 12'h000;
    rom[10648] = 12'h000;
    rom[10649] = 12'h000;
    rom[10650] = 12'h000;
    rom[10651] = 12'h000;
    rom[10652] = 12'h000;
    rom[10653] = 12'h000;
    rom[10654] = 12'h000;
    rom[10655] = 12'h000;
    rom[10656] = 12'h000;
    rom[10657] = 12'h000;
    rom[10658] = 12'h000;
    rom[10659] = 12'h000;
    rom[10660] = 12'h000;
    rom[10661] = 12'h000;
    rom[10662] = 12'h000;
    rom[10663] = 12'h000;
    rom[10664] = 12'h000;
    rom[10665] = 12'h000;
    rom[10666] = 12'h000;
    rom[10667] = 12'h000;
    rom[10668] = 12'h000;
    rom[10669] = 12'h000;
    rom[10670] = 12'h000;
    rom[10671] = 12'h000;
    rom[10672] = 12'h000;
    rom[10673] = 12'h000;
    rom[10674] = 12'h000;
    rom[10675] = 12'h000;
    rom[10676] = 12'h000;
    rom[10677] = 12'h000;
    rom[10678] = 12'h000;
    rom[10679] = 12'h000;
    rom[10680] = 12'h000;
    rom[10681] = 12'h000;
    rom[10682] = 12'h000;
    rom[10683] = 12'h000;
    rom[10684] = 12'h000;
    rom[10685] = 12'h000;
    rom[10686] = 12'h000;
    rom[10687] = 12'h000;
    rom[10688] = 12'h000;
    rom[10689] = 12'h000;
    rom[10690] = 12'h000;
    rom[10691] = 12'h000;
    rom[10692] = 12'h000;
    rom[10693] = 12'h000;
    rom[10694] = 12'h000;
    rom[10695] = 12'h000;
    rom[10696] = 12'h000;
    rom[10697] = 12'h000;
    rom[10698] = 12'h000;
    rom[10699] = 12'h000;
    rom[10700] = 12'h000;
    rom[10701] = 12'h000;
    rom[10702] = 12'h000;
    rom[10703] = 12'h000;
    rom[10704] = 12'h000;
    rom[10705] = 12'h000;
    rom[10706] = 12'h000;
    rom[10707] = 12'h000;
    rom[10708] = 12'h000;
    rom[10709] = 12'h000;
    rom[10710] = 12'h000;
    rom[10711] = 12'h000;
    rom[10712] = 12'h000;
    rom[10713] = 12'h000;
    rom[10714] = 12'h000;
    rom[10715] = 12'h000;
    rom[10716] = 12'h000;
    rom[10717] = 12'h000;
    rom[10718] = 12'h000;
    rom[10719] = 12'h000;
    rom[10720] = 12'h000;
    rom[10721] = 12'h000;
    rom[10722] = 12'h000;
    rom[10723] = 12'h000;
    rom[10724] = 12'h000;
    rom[10725] = 12'h000;
    rom[10726] = 12'h000;
    rom[10727] = 12'h000;
    rom[10728] = 12'h000;
    rom[10729] = 12'h000;
    rom[10730] = 12'h000;
    rom[10731] = 12'h000;
    rom[10732] = 12'h000;
    rom[10733] = 12'h3a2;
    rom[10734] = 12'h3a2;
    rom[10735] = 12'h3a2;
    rom[10736] = 12'h3a2;
    rom[10737] = 12'h3a2;
    rom[10738] = 12'h3a2;
    rom[10739] = 12'h3a2;
    rom[10740] = 12'h3a2;
    rom[10741] = 12'h3a2;
    rom[10742] = 12'h3a2;
    rom[10743] = 12'h3a2;
    rom[10744] = 12'h3a2;
    rom[10745] = 12'h3a2;
    rom[10746] = 12'h3a2;
    rom[10747] = 12'h3a2;
    rom[10748] = 12'h3a2;
    rom[10749] = 12'h000;
    rom[10750] = 12'h000;
    rom[10751] = 12'h000;
    rom[10752] = 12'h000;
    rom[10753] = 12'h000;
    rom[10754] = 12'h000;
    rom[10755] = 12'h2dc;
    rom[10756] = 12'h2dc;
    rom[10757] = 12'h2dc;
    rom[10758] = 12'h2dc;
    rom[10759] = 12'h2dc;
    rom[10760] = 12'h2dc;
    rom[10761] = 12'h2dd;
    rom[10762] = 12'h2dd;
    rom[10763] = 12'h2dd;
    rom[10764] = 12'h2dd;
    rom[10765] = 12'h2dd;
    rom[10766] = 12'h2dd;
    rom[10767] = 12'h2dd;
    rom[10768] = 12'h2dd;
    rom[10769] = 12'h2dd;
    rom[10770] = 12'h2dd;
    rom[10771] = 12'h000;
    rom[10772] = 12'h000;
    rom[10773] = 12'h000;
    rom[10774] = 12'h000;
    rom[10775] = 12'h000;
    rom[10776] = 12'h000;
    rom[10777] = 12'h000;
    rom[10778] = 12'h000;
    rom[10779] = 12'h000;
    rom[10780] = 12'h000;
    rom[10781] = 12'h000;
    rom[10782] = 12'h000;
    rom[10783] = 12'h000;
    rom[10784] = 12'h000;
    rom[10785] = 12'h000;
    rom[10786] = 12'h000;
    rom[10787] = 12'h000;
    rom[10788] = 12'h000;
    rom[10789] = 12'h000;
    rom[10790] = 12'h000;
    rom[10791] = 12'h000;
    rom[10792] = 12'h000;
    rom[10793] = 12'h000;
    rom[10794] = 12'h000;
    rom[10795] = 12'h000;
    rom[10796] = 12'h000;
    rom[10797] = 12'h000;
    rom[10798] = 12'h000;
    rom[10799] = 12'h000;
    rom[10800] = 12'h000;
    rom[10801] = 12'h000;
    rom[10802] = 12'h000;
    rom[10803] = 12'h000;
    rom[10804] = 12'h000;
    rom[10805] = 12'h000;
    rom[10806] = 12'h000;
    rom[10807] = 12'h000;
    rom[10808] = 12'h000;
    rom[10809] = 12'h000;
    rom[10810] = 12'h000;
    rom[10811] = 12'h000;
    rom[10812] = 12'h000;
    rom[10813] = 12'h000;
    rom[10814] = 12'h000;
    rom[10815] = 12'h000;
    rom[10816] = 12'h000;
    rom[10817] = 12'h000;
    rom[10818] = 12'h000;
    rom[10819] = 12'h000;
    rom[10820] = 12'h000;
    rom[10821] = 12'h000;
    rom[10822] = 12'h000;
    rom[10823] = 12'h000;
    rom[10824] = 12'h000;
    rom[10825] = 12'h000;
    rom[10826] = 12'h000;
    rom[10827] = 12'h000;
    rom[10828] = 12'h000;
    rom[10829] = 12'h000;
    rom[10830] = 12'h000;
    rom[10831] = 12'h000;
    rom[10832] = 12'h000;
    rom[10833] = 12'h000;
    rom[10834] = 12'h000;
    rom[10835] = 12'h000;
    rom[10836] = 12'h000;
    rom[10837] = 12'h000;
    rom[10838] = 12'h000;
    rom[10839] = 12'h000;
    rom[10840] = 12'h000;
    rom[10841] = 12'h000;
    rom[10842] = 12'h000;
    rom[10843] = 12'h000;
    rom[10844] = 12'h000;
    rom[10845] = 12'h000;
    rom[10846] = 12'h000;
    rom[10847] = 12'h000;
    rom[10848] = 12'h000;
    rom[10849] = 12'h000;
    rom[10850] = 12'h000;
    rom[10851] = 12'h000;
    rom[10852] = 12'h000;
    rom[10853] = 12'h000;
    rom[10854] = 12'h000;
    rom[10855] = 12'h000;
    rom[10856] = 12'h000;
    rom[10857] = 12'h000;
    rom[10858] = 12'h000;
    rom[10859] = 12'h000;
    rom[10860] = 12'h000;
    rom[10861] = 12'h3a2;
    rom[10862] = 12'h3a2;
    rom[10863] = 12'h3a2;
    rom[10864] = 12'h3a2;
    rom[10865] = 12'h3a2;
    rom[10866] = 12'h3a2;
    rom[10867] = 12'h3a2;
    rom[10868] = 12'h3a2;
    rom[10869] = 12'h3a2;
    rom[10870] = 12'h3a2;
    rom[10871] = 12'h3a2;
    rom[10872] = 12'h3a2;
    rom[10873] = 12'h3a2;
    rom[10874] = 12'h3a2;
    rom[10875] = 12'h3a2;
    rom[10876] = 12'h3a2;
    rom[10877] = 12'h000;
    rom[10878] = 12'h000;
    rom[10879] = 12'h000;
    rom[10880] = 12'h000;
    rom[10881] = 12'h000;
    rom[10882] = 12'h000;
    rom[10883] = 12'h000;
    rom[10884] = 12'h2dc;
    rom[10885] = 12'h2dc;
    rom[10886] = 12'h2dd;
    rom[10887] = 12'h2dd;
    rom[10888] = 12'h2dd;
    rom[10889] = 12'h2dd;
    rom[10890] = 12'h2dd;
    rom[10891] = 12'h2dd;
    rom[10892] = 12'h2dd;
    rom[10893] = 12'h2dd;
    rom[10894] = 12'h2dd;
    rom[10895] = 12'h2dd;
    rom[10896] = 12'h2ed;
    rom[10897] = 12'h1ed;
    rom[10898] = 12'h1ed;
    rom[10899] = 12'h1ed;
    rom[10900] = 12'h000;
    rom[10901] = 12'h000;
    rom[10902] = 12'h000;
    rom[10903] = 12'h000;
    rom[10904] = 12'h000;
    rom[10905] = 12'h000;
    rom[10906] = 12'h000;
    rom[10907] = 12'h000;
    rom[10908] = 12'h000;
    rom[10909] = 12'h000;
    rom[10910] = 12'h000;
    rom[10911] = 12'h000;
    rom[10912] = 12'h000;
    rom[10913] = 12'h000;
    rom[10914] = 12'h000;
    rom[10915] = 12'h000;
    rom[10916] = 12'h000;
    rom[10917] = 12'h000;
    rom[10918] = 12'h000;
    rom[10919] = 12'h000;
    rom[10920] = 12'h000;
    rom[10921] = 12'h000;
    rom[10922] = 12'h000;
    rom[10923] = 12'h000;
    rom[10924] = 12'h000;
    rom[10925] = 12'h000;
    rom[10926] = 12'h000;
    rom[10927] = 12'h000;
    rom[10928] = 12'h000;
    rom[10929] = 12'h000;
    rom[10930] = 12'h000;
    rom[10931] = 12'h000;
    rom[10932] = 12'h000;
    rom[10933] = 12'h000;
    rom[10934] = 12'h000;
    rom[10935] = 12'h000;
    rom[10936] = 12'h000;
    rom[10937] = 12'h000;
    rom[10938] = 12'h000;
    rom[10939] = 12'h000;
    rom[10940] = 12'h000;
    rom[10941] = 12'h000;
    rom[10942] = 12'h000;
    rom[10943] = 12'h000;
    rom[10944] = 12'h000;
    rom[10945] = 12'h000;
    rom[10946] = 12'h000;
    rom[10947] = 12'h000;
    rom[10948] = 12'h000;
    rom[10949] = 12'h000;
    rom[10950] = 12'h000;
    rom[10951] = 12'h000;
    rom[10952] = 12'h000;
    rom[10953] = 12'h000;
    rom[10954] = 12'h000;
    rom[10955] = 12'h000;
    rom[10956] = 12'h000;
    rom[10957] = 12'h000;
    rom[10958] = 12'h000;
    rom[10959] = 12'h000;
    rom[10960] = 12'h000;
    rom[10961] = 12'h000;
    rom[10962] = 12'h000;
    rom[10963] = 12'h000;
    rom[10964] = 12'h000;
    rom[10965] = 12'h000;
    rom[10966] = 12'h000;
    rom[10967] = 12'h000;
    rom[10968] = 12'h000;
    rom[10969] = 12'h000;
    rom[10970] = 12'h000;
    rom[10971] = 12'h000;
    rom[10972] = 12'h000;
    rom[10973] = 12'h000;
    rom[10974] = 12'h000;
    rom[10975] = 12'h000;
    rom[10976] = 12'h000;
    rom[10977] = 12'h000;
    rom[10978] = 12'h000;
    rom[10979] = 12'h000;
    rom[10980] = 12'h000;
    rom[10981] = 12'h000;
    rom[10982] = 12'h000;
    rom[10983] = 12'h000;
    rom[10984] = 12'h000;
    rom[10985] = 12'h000;
    rom[10986] = 12'h000;
    rom[10987] = 12'h000;
    rom[10988] = 12'h3a2;
    rom[10989] = 12'h3a2;
    rom[10990] = 12'h3a2;
    rom[10991] = 12'h3a2;
    rom[10992] = 12'h3a2;
    rom[10993] = 12'h3a2;
    rom[10994] = 12'h3a2;
    rom[10995] = 12'h3a2;
    rom[10996] = 12'h3a2;
    rom[10997] = 12'h3a2;
    rom[10998] = 12'h3a2;
    rom[10999] = 12'h3a2;
    rom[11000] = 12'h3a2;
    rom[11001] = 12'h3a2;
    rom[11002] = 12'h3a2;
    rom[11003] = 12'h3a2;
    rom[11004] = 12'h000;
    rom[11005] = 12'h000;
    rom[11006] = 12'h000;
    rom[11007] = 12'h000;
    rom[11008] = 12'h000;
    rom[11009] = 12'h000;
    rom[11010] = 12'h000;
    rom[11011] = 12'h000;
    rom[11012] = 12'h2dd;
    rom[11013] = 12'h2dd;
    rom[11014] = 12'h2dd;
    rom[11015] = 12'h2dd;
    rom[11016] = 12'h2dd;
    rom[11017] = 12'h2dd;
    rom[11018] = 12'h2dd;
    rom[11019] = 12'h2dd;
    rom[11020] = 12'h2dd;
    rom[11021] = 12'h2dd;
    rom[11022] = 12'h1ed;
    rom[11023] = 12'h1ed;
    rom[11024] = 12'h1ed;
    rom[11025] = 12'h1ed;
    rom[11026] = 12'h1ed;
    rom[11027] = 12'h1ed;
    rom[11028] = 12'h000;
    rom[11029] = 12'h000;
    rom[11030] = 12'h000;
    rom[11031] = 12'h000;
    rom[11032] = 12'h000;
    rom[11033] = 12'h000;
    rom[11034] = 12'h000;
    rom[11035] = 12'h000;
    rom[11036] = 12'h000;
    rom[11037] = 12'h000;
    rom[11038] = 12'h000;
    rom[11039] = 12'h000;
    rom[11040] = 12'h000;
    rom[11041] = 12'h000;
    rom[11042] = 12'h000;
    rom[11043] = 12'h000;
    rom[11044] = 12'h000;
    rom[11045] = 12'h000;
    rom[11046] = 12'h000;
    rom[11047] = 12'h000;
    rom[11048] = 12'h000;
    rom[11049] = 12'h000;
    rom[11050] = 12'h000;
    rom[11051] = 12'h000;
    rom[11052] = 12'h000;
    rom[11053] = 12'h000;
    rom[11054] = 12'h000;
    rom[11055] = 12'h000;
    rom[11056] = 12'h000;
    rom[11057] = 12'h000;
    rom[11058] = 12'h000;
    rom[11059] = 12'h000;
    rom[11060] = 12'h000;
    rom[11061] = 12'h000;
    rom[11062] = 12'h000;
    rom[11063] = 12'h000;
    rom[11064] = 12'h000;
    rom[11065] = 12'h000;
    rom[11066] = 12'h000;
    rom[11067] = 12'h000;
    rom[11068] = 12'h000;
    rom[11069] = 12'h000;
    rom[11070] = 12'h000;
    rom[11071] = 12'h000;
    rom[11072] = 12'h000;
    rom[11073] = 12'h000;
    rom[11074] = 12'h000;
    rom[11075] = 12'h000;
    rom[11076] = 12'h000;
    rom[11077] = 12'h000;
    rom[11078] = 12'h000;
    rom[11079] = 12'h000;
    rom[11080] = 12'h000;
    rom[11081] = 12'h000;
    rom[11082] = 12'h000;
    rom[11083] = 12'h000;
    rom[11084] = 12'h000;
    rom[11085] = 12'h000;
    rom[11086] = 12'h000;
    rom[11087] = 12'h000;
    rom[11088] = 12'h000;
    rom[11089] = 12'h000;
    rom[11090] = 12'h000;
    rom[11091] = 12'h000;
    rom[11092] = 12'h000;
    rom[11093] = 12'h000;
    rom[11094] = 12'h000;
    rom[11095] = 12'h000;
    rom[11096] = 12'h000;
    rom[11097] = 12'h000;
    rom[11098] = 12'h000;
    rom[11099] = 12'h000;
    rom[11100] = 12'h000;
    rom[11101] = 12'h000;
    rom[11102] = 12'h000;
    rom[11103] = 12'h000;
    rom[11104] = 12'h000;
    rom[11105] = 12'h000;
    rom[11106] = 12'h000;
    rom[11107] = 12'h000;
    rom[11108] = 12'h000;
    rom[11109] = 12'h000;
    rom[11110] = 12'h000;
    rom[11111] = 12'h000;
    rom[11112] = 12'h000;
    rom[11113] = 12'h000;
    rom[11114] = 12'h000;
    rom[11115] = 12'h000;
    rom[11116] = 12'h3a2;
    rom[11117] = 12'h3a2;
    rom[11118] = 12'h3a2;
    rom[11119] = 12'h3a2;
    rom[11120] = 12'h3a2;
    rom[11121] = 12'h3a2;
    rom[11122] = 12'h3a2;
    rom[11123] = 12'h3a2;
    rom[11124] = 12'h3a2;
    rom[11125] = 12'h3a2;
    rom[11126] = 12'h3a2;
    rom[11127] = 12'h3a2;
    rom[11128] = 12'h3a2;
    rom[11129] = 12'h3a2;
    rom[11130] = 12'h3a2;
    rom[11131] = 12'h3a2;
    rom[11132] = 12'h000;
    rom[11133] = 12'h000;
    rom[11134] = 12'h000;
    rom[11135] = 12'h000;
    rom[11136] = 12'h000;
    rom[11137] = 12'h000;
    rom[11138] = 12'h000;
    rom[11139] = 12'h000;
    rom[11140] = 12'h2dd;
    rom[11141] = 12'h2dd;
    rom[11142] = 12'h2dd;
    rom[11143] = 12'h2dd;
    rom[11144] = 12'h2dd;
    rom[11145] = 12'h2dd;
    rom[11146] = 12'h2dd;
    rom[11147] = 12'h1ed;
    rom[11148] = 12'h1ed;
    rom[11149] = 12'h1ed;
    rom[11150] = 12'h1ed;
    rom[11151] = 12'h1ed;
    rom[11152] = 12'h1ed;
    rom[11153] = 12'h1ed;
    rom[11154] = 12'h1ed;
    rom[11155] = 12'h1ed;
    rom[11156] = 12'h1ed;
    rom[11157] = 12'h000;
    rom[11158] = 12'h000;
    rom[11159] = 12'h000;
    rom[11160] = 12'h000;
    rom[11161] = 12'h000;
    rom[11162] = 12'h000;
    rom[11163] = 12'h000;
    rom[11164] = 12'h000;
    rom[11165] = 12'h000;
    rom[11166] = 12'h000;
    rom[11167] = 12'h000;
    rom[11168] = 12'h000;
    rom[11169] = 12'h000;
    rom[11170] = 12'h000;
    rom[11171] = 12'h000;
    rom[11172] = 12'h000;
    rom[11173] = 12'h000;
    rom[11174] = 12'h000;
    rom[11175] = 12'h000;
    rom[11176] = 12'h000;
    rom[11177] = 12'h000;
    rom[11178] = 12'h000;
    rom[11179] = 12'h000;
    rom[11180] = 12'h000;
    rom[11181] = 12'h000;
    rom[11182] = 12'h000;
    rom[11183] = 12'h000;
    rom[11184] = 12'h000;
    rom[11185] = 12'h000;
    rom[11186] = 12'h000;
    rom[11187] = 12'h000;
    rom[11188] = 12'h000;
    rom[11189] = 12'h000;
    rom[11190] = 12'h000;
    rom[11191] = 12'h000;
    rom[11192] = 12'h000;
    rom[11193] = 12'h000;
    rom[11194] = 12'h000;
    rom[11195] = 12'h000;
    rom[11196] = 12'h000;
    rom[11197] = 12'h000;
    rom[11198] = 12'h000;
    rom[11199] = 12'h000;
    rom[11200] = 12'h000;
    rom[11201] = 12'h000;
    rom[11202] = 12'h000;
    rom[11203] = 12'h000;
    rom[11204] = 12'h000;
    rom[11205] = 12'h000;
    rom[11206] = 12'h000;
    rom[11207] = 12'h000;
    rom[11208] = 12'h000;
    rom[11209] = 12'h000;
    rom[11210] = 12'h000;
    rom[11211] = 12'h000;
    rom[11212] = 12'h000;
    rom[11213] = 12'h000;
    rom[11214] = 12'h000;
    rom[11215] = 12'h000;
    rom[11216] = 12'h000;
    rom[11217] = 12'h000;
    rom[11218] = 12'h000;
    rom[11219] = 12'h000;
    rom[11220] = 12'h000;
    rom[11221] = 12'h000;
    rom[11222] = 12'h000;
    rom[11223] = 12'h000;
    rom[11224] = 12'h000;
    rom[11225] = 12'h000;
    rom[11226] = 12'h000;
    rom[11227] = 12'h000;
    rom[11228] = 12'h000;
    rom[11229] = 12'h000;
    rom[11230] = 12'h000;
    rom[11231] = 12'h000;
    rom[11232] = 12'h000;
    rom[11233] = 12'h000;
    rom[11234] = 12'h000;
    rom[11235] = 12'h000;
    rom[11236] = 12'h000;
    rom[11237] = 12'h000;
    rom[11238] = 12'h000;
    rom[11239] = 12'h000;
    rom[11240] = 12'h000;
    rom[11241] = 12'h000;
    rom[11242] = 12'h000;
    rom[11243] = 12'h3a2;
    rom[11244] = 12'h3a2;
    rom[11245] = 12'h3a2;
    rom[11246] = 12'h3a2;
    rom[11247] = 12'h3a2;
    rom[11248] = 12'h3a2;
    rom[11249] = 12'h3a2;
    rom[11250] = 12'h3a2;
    rom[11251] = 12'h3a2;
    rom[11252] = 12'h3a2;
    rom[11253] = 12'h3a2;
    rom[11254] = 12'h3a2;
    rom[11255] = 12'h3a2;
    rom[11256] = 12'h3a2;
    rom[11257] = 12'h3a2;
    rom[11258] = 12'h3a2;
    rom[11259] = 12'h3a2;
    rom[11260] = 12'h000;
    rom[11261] = 12'h000;
    rom[11262] = 12'h000;
    rom[11263] = 12'h000;
    rom[11264] = 12'h000;
    rom[11265] = 12'h000;
    rom[11266] = 12'h000;
    rom[11267] = 12'h000;
    rom[11268] = 12'h000;
    rom[11269] = 12'h2dd;
    rom[11270] = 12'h2dd;
    rom[11271] = 12'h2dd;
    rom[11272] = 12'h1ed;
    rom[11273] = 12'h1ed;
    rom[11274] = 12'h1ed;
    rom[11275] = 12'h1ed;
    rom[11276] = 12'h1ed;
    rom[11277] = 12'h1ed;
    rom[11278] = 12'h1ed;
    rom[11279] = 12'h1ed;
    rom[11280] = 12'h1ed;
    rom[11281] = 12'h1ed;
    rom[11282] = 12'h1ed;
    rom[11283] = 12'h1ee;
    rom[11284] = 12'h1ee;
    rom[11285] = 12'h000;
    rom[11286] = 12'h000;
    rom[11287] = 12'h000;
    rom[11288] = 12'h000;
    rom[11289] = 12'h000;
    rom[11290] = 12'h000;
    rom[11291] = 12'h000;
    rom[11292] = 12'h000;
    rom[11293] = 12'h000;
    rom[11294] = 12'h000;
    rom[11295] = 12'h000;
    rom[11296] = 12'h000;
    rom[11297] = 12'h000;
    rom[11298] = 12'h000;
    rom[11299] = 12'h000;
    rom[11300] = 12'h000;
    rom[11301] = 12'h000;
    rom[11302] = 12'h000;
    rom[11303] = 12'h000;
    rom[11304] = 12'h000;
    rom[11305] = 12'h000;
    rom[11306] = 12'h000;
    rom[11307] = 12'h000;
    rom[11308] = 12'h000;
    rom[11309] = 12'h000;
    rom[11310] = 12'h000;
    rom[11311] = 12'h000;
    rom[11312] = 12'h000;
    rom[11313] = 12'h000;
    rom[11314] = 12'h000;
    rom[11315] = 12'h000;
    rom[11316] = 12'h000;
    rom[11317] = 12'h000;
    rom[11318] = 12'h000;
    rom[11319] = 12'h000;
    rom[11320] = 12'h000;
    rom[11321] = 12'h000;
    rom[11322] = 12'h000;
    rom[11323] = 12'h000;
    rom[11324] = 12'h000;
    rom[11325] = 12'h000;
    rom[11326] = 12'h000;
    rom[11327] = 12'h000;
    rom[11328] = 12'h000;
    rom[11329] = 12'h000;
    rom[11330] = 12'h000;
    rom[11331] = 12'h000;
    rom[11332] = 12'h000;
    rom[11333] = 12'h000;
    rom[11334] = 12'h000;
    rom[11335] = 12'h000;
    rom[11336] = 12'h000;
    rom[11337] = 12'h000;
    rom[11338] = 12'h000;
    rom[11339] = 12'h000;
    rom[11340] = 12'h000;
    rom[11341] = 12'h000;
    rom[11342] = 12'h000;
    rom[11343] = 12'h000;
    rom[11344] = 12'h000;
    rom[11345] = 12'h000;
    rom[11346] = 12'h000;
    rom[11347] = 12'h000;
    rom[11348] = 12'h000;
    rom[11349] = 12'h000;
    rom[11350] = 12'h000;
    rom[11351] = 12'h000;
    rom[11352] = 12'h000;
    rom[11353] = 12'h000;
    rom[11354] = 12'h000;
    rom[11355] = 12'h000;
    rom[11356] = 12'h000;
    rom[11357] = 12'h000;
    rom[11358] = 12'h000;
    rom[11359] = 12'h000;
    rom[11360] = 12'h000;
    rom[11361] = 12'h000;
    rom[11362] = 12'h000;
    rom[11363] = 12'h000;
    rom[11364] = 12'h000;
    rom[11365] = 12'h000;
    rom[11366] = 12'h000;
    rom[11367] = 12'h000;
    rom[11368] = 12'h000;
    rom[11369] = 12'h000;
    rom[11370] = 12'h000;
    rom[11371] = 12'h3a2;
    rom[11372] = 12'h3a2;
    rom[11373] = 12'h3a2;
    rom[11374] = 12'h3a2;
    rom[11375] = 12'h3a2;
    rom[11376] = 12'h3a2;
    rom[11377] = 12'h3a2;
    rom[11378] = 12'h3a2;
    rom[11379] = 12'h3a2;
    rom[11380] = 12'h3a2;
    rom[11381] = 12'h3a2;
    rom[11382] = 12'h3a2;
    rom[11383] = 12'h3a2;
    rom[11384] = 12'h3a2;
    rom[11385] = 12'h3a2;
    rom[11386] = 12'h3a2;
    rom[11387] = 12'h000;
    rom[11388] = 12'h000;
    rom[11389] = 12'h000;
    rom[11390] = 12'h000;
    rom[11391] = 12'h000;
    rom[11392] = 12'h000;
    rom[11393] = 12'h000;
    rom[11394] = 12'h000;
    rom[11395] = 12'h000;
    rom[11396] = 12'h000;
    rom[11397] = 12'h1ed;
    rom[11398] = 12'h1ed;
    rom[11399] = 12'h1ed;
    rom[11400] = 12'h1ed;
    rom[11401] = 12'h1ed;
    rom[11402] = 12'h1ed;
    rom[11403] = 12'h1ed;
    rom[11404] = 12'h1ed;
    rom[11405] = 12'h1ed;
    rom[11406] = 12'h1ed;
    rom[11407] = 12'h1ed;
    rom[11408] = 12'h1ee;
    rom[11409] = 12'h1ee;
    rom[11410] = 12'h1ee;
    rom[11411] = 12'h1ee;
    rom[11412] = 12'h1ee;
    rom[11413] = 12'h1ee;
    rom[11414] = 12'h000;
    rom[11415] = 12'h000;
    rom[11416] = 12'h000;
    rom[11417] = 12'h000;
    rom[11418] = 12'h000;
    rom[11419] = 12'h000;
    rom[11420] = 12'h000;
    rom[11421] = 12'h000;
    rom[11422] = 12'h000;
    rom[11423] = 12'h000;
    rom[11424] = 12'h000;
    rom[11425] = 12'h000;
    rom[11426] = 12'h000;
    rom[11427] = 12'h000;
    rom[11428] = 12'h000;
    rom[11429] = 12'h000;
    rom[11430] = 12'h000;
    rom[11431] = 12'h000;
    rom[11432] = 12'h000;
    rom[11433] = 12'h000;
    rom[11434] = 12'h000;
    rom[11435] = 12'h000;
    rom[11436] = 12'h000;
    rom[11437] = 12'h000;
    rom[11438] = 12'h000;
    rom[11439] = 12'h000;
    rom[11440] = 12'h000;
    rom[11441] = 12'h000;
    rom[11442] = 12'h000;
    rom[11443] = 12'h000;
    rom[11444] = 12'h000;
    rom[11445] = 12'h000;
    rom[11446] = 12'h000;
    rom[11447] = 12'h000;
    rom[11448] = 12'h000;
    rom[11449] = 12'h000;
    rom[11450] = 12'h000;
    rom[11451] = 12'h000;
    rom[11452] = 12'h000;
    rom[11453] = 12'h000;
    rom[11454] = 12'h000;
    rom[11455] = 12'h000;
    rom[11456] = 12'h000;
    rom[11457] = 12'h000;
    rom[11458] = 12'h000;
    rom[11459] = 12'h000;
    rom[11460] = 12'h000;
    rom[11461] = 12'h000;
    rom[11462] = 12'h000;
    rom[11463] = 12'h000;
    rom[11464] = 12'h000;
    rom[11465] = 12'h000;
    rom[11466] = 12'h000;
    rom[11467] = 12'h000;
    rom[11468] = 12'h000;
    rom[11469] = 12'h000;
    rom[11470] = 12'h000;
    rom[11471] = 12'h000;
    rom[11472] = 12'h000;
    rom[11473] = 12'h000;
    rom[11474] = 12'h000;
    rom[11475] = 12'h000;
    rom[11476] = 12'h000;
    rom[11477] = 12'h000;
    rom[11478] = 12'h000;
    rom[11479] = 12'h000;
    rom[11480] = 12'h000;
    rom[11481] = 12'h000;
    rom[11482] = 12'h000;
    rom[11483] = 12'h000;
    rom[11484] = 12'h000;
    rom[11485] = 12'h000;
    rom[11486] = 12'h000;
    rom[11487] = 12'h000;
    rom[11488] = 12'h000;
    rom[11489] = 12'h000;
    rom[11490] = 12'h000;
    rom[11491] = 12'h000;
    rom[11492] = 12'h000;
    rom[11493] = 12'h000;
    rom[11494] = 12'h000;
    rom[11495] = 12'h000;
    rom[11496] = 12'h000;
    rom[11497] = 12'h000;
    rom[11498] = 12'h3a2;
    rom[11499] = 12'h3a2;
    rom[11500] = 12'h3a2;
    rom[11501] = 12'h3a2;
    rom[11502] = 12'h3a2;
    rom[11503] = 12'h3a2;
    rom[11504] = 12'h3a2;
    rom[11505] = 12'h3a2;
    rom[11506] = 12'h3a2;
    rom[11507] = 12'h3a2;
    rom[11508] = 12'h3a2;
    rom[11509] = 12'h3a2;
    rom[11510] = 12'h3a2;
    rom[11511] = 12'h3a2;
    rom[11512] = 12'h3a2;
    rom[11513] = 12'h3a2;
    rom[11514] = 12'h3a2;
    rom[11515] = 12'h000;
    rom[11516] = 12'h000;
    rom[11517] = 12'h000;
    rom[11518] = 12'h000;
    rom[11519] = 12'h000;
    rom[11520] = 12'h000;
    rom[11521] = 12'h000;
    rom[11522] = 12'h000;
    rom[11523] = 12'h000;
    rom[11524] = 12'h000;
    rom[11525] = 12'h000;
    rom[11526] = 12'h1ed;
    rom[11527] = 12'h1ed;
    rom[11528] = 12'h1ed;
    rom[11529] = 12'h1ed;
    rom[11530] = 12'h1ed;
    rom[11531] = 12'h1ed;
    rom[11532] = 12'h1ed;
    rom[11533] = 12'h1ee;
    rom[11534] = 12'h1ee;
    rom[11535] = 12'h1ee;
    rom[11536] = 12'h1ee;
    rom[11537] = 12'h1ee;
    rom[11538] = 12'h1ee;
    rom[11539] = 12'h1ee;
    rom[11540] = 12'h1ee;
    rom[11541] = 12'h1ee;
    rom[11542] = 12'h1ee;
    rom[11543] = 12'h000;
    rom[11544] = 12'h000;
    rom[11545] = 12'h000;
    rom[11546] = 12'h000;
    rom[11547] = 12'h000;
    rom[11548] = 12'h000;
    rom[11549] = 12'h000;
    rom[11550] = 12'h000;
    rom[11551] = 12'h000;
    rom[11552] = 12'h000;
    rom[11553] = 12'h000;
    rom[11554] = 12'h000;
    rom[11555] = 12'h000;
    rom[11556] = 12'h000;
    rom[11557] = 12'h000;
    rom[11558] = 12'h000;
    rom[11559] = 12'h000;
    rom[11560] = 12'h000;
    rom[11561] = 12'h000;
    rom[11562] = 12'h000;
    rom[11563] = 12'h000;
    rom[11564] = 12'h000;
    rom[11565] = 12'h000;
    rom[11566] = 12'h000;
    rom[11567] = 12'h000;
    rom[11568] = 12'h000;
    rom[11569] = 12'h000;
    rom[11570] = 12'h000;
    rom[11571] = 12'h000;
    rom[11572] = 12'h000;
    rom[11573] = 12'h000;
    rom[11574] = 12'h000;
    rom[11575] = 12'h000;
    rom[11576] = 12'h000;
    rom[11577] = 12'h000;
    rom[11578] = 12'h000;
    rom[11579] = 12'h000;
    rom[11580] = 12'h000;
    rom[11581] = 12'h000;
    rom[11582] = 12'h000;
    rom[11583] = 12'h000;
    rom[11584] = 12'h000;
    rom[11585] = 12'h000;
    rom[11586] = 12'h000;
    rom[11587] = 12'h000;
    rom[11588] = 12'h000;
    rom[11589] = 12'h000;
    rom[11590] = 12'h000;
    rom[11591] = 12'h000;
    rom[11592] = 12'h000;
    rom[11593] = 12'h000;
    rom[11594] = 12'h000;
    rom[11595] = 12'h000;
    rom[11596] = 12'h000;
    rom[11597] = 12'h000;
    rom[11598] = 12'h000;
    rom[11599] = 12'h000;
    rom[11600] = 12'h000;
    rom[11601] = 12'h000;
    rom[11602] = 12'h000;
    rom[11603] = 12'h000;
    rom[11604] = 12'h000;
    rom[11605] = 12'h000;
    rom[11606] = 12'h000;
    rom[11607] = 12'h000;
    rom[11608] = 12'h000;
    rom[11609] = 12'h000;
    rom[11610] = 12'h000;
    rom[11611] = 12'h000;
    rom[11612] = 12'h000;
    rom[11613] = 12'h000;
    rom[11614] = 12'h000;
    rom[11615] = 12'h000;
    rom[11616] = 12'h000;
    rom[11617] = 12'h000;
    rom[11618] = 12'h000;
    rom[11619] = 12'h000;
    rom[11620] = 12'h000;
    rom[11621] = 12'h000;
    rom[11622] = 12'h000;
    rom[11623] = 12'h000;
    rom[11624] = 12'h000;
    rom[11625] = 12'h392;
    rom[11626] = 12'h3a2;
    rom[11627] = 12'h3a2;
    rom[11628] = 12'h3a2;
    rom[11629] = 12'h3a2;
    rom[11630] = 12'h3a2;
    rom[11631] = 12'h3a2;
    rom[11632] = 12'h3a2;
    rom[11633] = 12'h3a2;
    rom[11634] = 12'h3a2;
    rom[11635] = 12'h3a2;
    rom[11636] = 12'h3a2;
    rom[11637] = 12'h3a2;
    rom[11638] = 12'h3a2;
    rom[11639] = 12'h3a2;
    rom[11640] = 12'h3a2;
    rom[11641] = 12'h3a2;
    rom[11642] = 12'h000;
    rom[11643] = 12'h000;
    rom[11644] = 12'h000;
    rom[11645] = 12'h000;
    rom[11646] = 12'h000;
    rom[11647] = 12'h000;
    rom[11648] = 12'h000;
    rom[11649] = 12'h000;
    rom[11650] = 12'h000;
    rom[11651] = 12'h000;
    rom[11652] = 12'h000;
    rom[11653] = 12'h000;
    rom[11654] = 12'h1ed;
    rom[11655] = 12'h1ed;
    rom[11656] = 12'h1ed;
    rom[11657] = 12'h1ed;
    rom[11658] = 12'h1ed;
    rom[11659] = 12'h1ee;
    rom[11660] = 12'h1ee;
    rom[11661] = 12'h1ee;
    rom[11662] = 12'h1ee;
    rom[11663] = 12'h1ee;
    rom[11664] = 12'h1ee;
    rom[11665] = 12'h1ee;
    rom[11666] = 12'h1ee;
    rom[11667] = 12'h1ee;
    rom[11668] = 12'h1ee;
    rom[11669] = 12'h1ee;
    rom[11670] = 12'h1ee;
    rom[11671] = 12'h000;
    rom[11672] = 12'h000;
    rom[11673] = 12'h000;
    rom[11674] = 12'h000;
    rom[11675] = 12'h000;
    rom[11676] = 12'h000;
    rom[11677] = 12'h000;
    rom[11678] = 12'h000;
    rom[11679] = 12'h000;
    rom[11680] = 12'h000;
    rom[11681] = 12'h000;
    rom[11682] = 12'h000;
    rom[11683] = 12'h000;
    rom[11684] = 12'h000;
    rom[11685] = 12'h000;
    rom[11686] = 12'h000;
    rom[11687] = 12'h000;
    rom[11688] = 12'h000;
    rom[11689] = 12'h000;
    rom[11690] = 12'h000;
    rom[11691] = 12'h000;
    rom[11692] = 12'h000;
    rom[11693] = 12'h000;
    rom[11694] = 12'h000;
    rom[11695] = 12'h000;
    rom[11696] = 12'h000;
    rom[11697] = 12'h000;
    rom[11698] = 12'h000;
    rom[11699] = 12'h000;
    rom[11700] = 12'h000;
    rom[11701] = 12'h000;
    rom[11702] = 12'h000;
    rom[11703] = 12'h000;
    rom[11704] = 12'h000;
    rom[11705] = 12'h000;
    rom[11706] = 12'h000;
    rom[11707] = 12'h000;
    rom[11708] = 12'h000;
    rom[11709] = 12'h000;
    rom[11710] = 12'h000;
    rom[11711] = 12'h000;
    rom[11712] = 12'h000;
    rom[11713] = 12'h000;
    rom[11714] = 12'h000;
    rom[11715] = 12'h000;
    rom[11716] = 12'h000;
    rom[11717] = 12'h000;
    rom[11718] = 12'h000;
    rom[11719] = 12'h000;
    rom[11720] = 12'h000;
    rom[11721] = 12'h000;
    rom[11722] = 12'h000;
    rom[11723] = 12'h000;
    rom[11724] = 12'h000;
    rom[11725] = 12'h000;
    rom[11726] = 12'h000;
    rom[11727] = 12'h000;
    rom[11728] = 12'h000;
    rom[11729] = 12'h000;
    rom[11730] = 12'h000;
    rom[11731] = 12'h000;
    rom[11732] = 12'h000;
    rom[11733] = 12'h000;
    rom[11734] = 12'h000;
    rom[11735] = 12'h000;
    rom[11736] = 12'h000;
    rom[11737] = 12'h000;
    rom[11738] = 12'h000;
    rom[11739] = 12'h000;
    rom[11740] = 12'h000;
    rom[11741] = 12'h000;
    rom[11742] = 12'h000;
    rom[11743] = 12'h000;
    rom[11744] = 12'h000;
    rom[11745] = 12'h000;
    rom[11746] = 12'h000;
    rom[11747] = 12'h000;
    rom[11748] = 12'h000;
    rom[11749] = 12'h000;
    rom[11750] = 12'h000;
    rom[11751] = 12'h000;
    rom[11752] = 12'h000;
    rom[11753] = 12'h3a2;
    rom[11754] = 12'h3a2;
    rom[11755] = 12'h3a2;
    rom[11756] = 12'h3a2;
    rom[11757] = 12'h3a2;
    rom[11758] = 12'h3a2;
    rom[11759] = 12'h3a2;
    rom[11760] = 12'h3a2;
    rom[11761] = 12'h3a2;
    rom[11762] = 12'h3a2;
    rom[11763] = 12'h3a2;
    rom[11764] = 12'h3a2;
    rom[11765] = 12'h3a2;
    rom[11766] = 12'h3a2;
    rom[11767] = 12'h3a2;
    rom[11768] = 12'h3a2;
    rom[11769] = 12'h3a2;
    rom[11770] = 12'h000;
    rom[11771] = 12'h000;
    rom[11772] = 12'h000;
    rom[11773] = 12'h000;
    rom[11774] = 12'h000;
    rom[11775] = 12'h000;
    rom[11776] = 12'h000;
    rom[11777] = 12'h000;
    rom[11778] = 12'h000;
    rom[11779] = 12'h000;
    rom[11780] = 12'h000;
    rom[11781] = 12'h000;
    rom[11782] = 12'h000;
    rom[11783] = 12'h1ed;
    rom[11784] = 12'h1ee;
    rom[11785] = 12'h1ee;
    rom[11786] = 12'h1ee;
    rom[11787] = 12'h1ee;
    rom[11788] = 12'h1ee;
    rom[11789] = 12'h1ee;
    rom[11790] = 12'h1ee;
    rom[11791] = 12'h1ee;
    rom[11792] = 12'h1ee;
    rom[11793] = 12'h1ee;
    rom[11794] = 12'h1ee;
    rom[11795] = 12'h1ee;
    rom[11796] = 12'h1ee;
    rom[11797] = 12'h1ee;
    rom[11798] = 12'h1ee;
    rom[11799] = 12'h1ee;
    rom[11800] = 12'h000;
    rom[11801] = 12'h000;
    rom[11802] = 12'h000;
    rom[11803] = 12'h000;
    rom[11804] = 12'h000;
    rom[11805] = 12'h000;
    rom[11806] = 12'h000;
    rom[11807] = 12'h000;
    rom[11808] = 12'h000;
    rom[11809] = 12'h000;
    rom[11810] = 12'h000;
    rom[11811] = 12'h000;
    rom[11812] = 12'h000;
    rom[11813] = 12'h000;
    rom[11814] = 12'h000;
    rom[11815] = 12'h000;
    rom[11816] = 12'h000;
    rom[11817] = 12'h000;
    rom[11818] = 12'h000;
    rom[11819] = 12'h000;
    rom[11820] = 12'h000;
    rom[11821] = 12'h000;
    rom[11822] = 12'h000;
    rom[11823] = 12'h000;
    rom[11824] = 12'h000;
    rom[11825] = 12'h000;
    rom[11826] = 12'h000;
    rom[11827] = 12'h000;
    rom[11828] = 12'h000;
    rom[11829] = 12'h000;
    rom[11830] = 12'h000;
    rom[11831] = 12'h000;
    rom[11832] = 12'h000;
    rom[11833] = 12'h000;
    rom[11834] = 12'h000;
    rom[11835] = 12'h000;
    rom[11836] = 12'h000;
    rom[11837] = 12'h000;
    rom[11838] = 12'h000;
    rom[11839] = 12'h000;
    rom[11840] = 12'h000;
    rom[11841] = 12'h000;
    rom[11842] = 12'h000;
    rom[11843] = 12'h000;
    rom[11844] = 12'h000;
    rom[11845] = 12'h000;
    rom[11846] = 12'h000;
    rom[11847] = 12'h000;
    rom[11848] = 12'h000;
    rom[11849] = 12'h000;
    rom[11850] = 12'h000;
    rom[11851] = 12'h000;
    rom[11852] = 12'h000;
    rom[11853] = 12'h000;
    rom[11854] = 12'h000;
    rom[11855] = 12'h000;
    rom[11856] = 12'h000;
    rom[11857] = 12'h000;
    rom[11858] = 12'h000;
    rom[11859] = 12'h000;
    rom[11860] = 12'h000;
    rom[11861] = 12'h000;
    rom[11862] = 12'h000;
    rom[11863] = 12'h000;
    rom[11864] = 12'h000;
    rom[11865] = 12'h000;
    rom[11866] = 12'h000;
    rom[11867] = 12'h000;
    rom[11868] = 12'h000;
    rom[11869] = 12'h000;
    rom[11870] = 12'h000;
    rom[11871] = 12'h000;
    rom[11872] = 12'h000;
    rom[11873] = 12'h000;
    rom[11874] = 12'h000;
    rom[11875] = 12'h000;
    rom[11876] = 12'h000;
    rom[11877] = 12'h000;
    rom[11878] = 12'h000;
    rom[11879] = 12'h000;
    rom[11880] = 12'h3a2;
    rom[11881] = 12'h3a2;
    rom[11882] = 12'h3a2;
    rom[11883] = 12'h3a2;
    rom[11884] = 12'h3a2;
    rom[11885] = 12'h3a2;
    rom[11886] = 12'h3a2;
    rom[11887] = 12'h3a2;
    rom[11888] = 12'h3a2;
    rom[11889] = 12'h3a2;
    rom[11890] = 12'h3a2;
    rom[11891] = 12'h3a2;
    rom[11892] = 12'h3a2;
    rom[11893] = 12'h3a2;
    rom[11894] = 12'h3a2;
    rom[11895] = 12'h3a2;
    rom[11896] = 12'h3a2;
    rom[11897] = 12'h000;
    rom[11898] = 12'h000;
    rom[11899] = 12'h000;
    rom[11900] = 12'h000;
    rom[11901] = 12'h000;
    rom[11902] = 12'h000;
    rom[11903] = 12'h000;
    rom[11904] = 12'h000;
    rom[11905] = 12'h000;
    rom[11906] = 12'h000;
    rom[11907] = 12'h000;
    rom[11908] = 12'h000;
    rom[11909] = 12'h000;
    rom[11910] = 12'h000;
    rom[11911] = 12'h1ee;
    rom[11912] = 12'h1ee;
    rom[11913] = 12'h1ee;
    rom[11914] = 12'h1ee;
    rom[11915] = 12'h1ee;
    rom[11916] = 12'h1ee;
    rom[11917] = 12'h1ee;
    rom[11918] = 12'h1ee;
    rom[11919] = 12'h1ee;
    rom[11920] = 12'h1ee;
    rom[11921] = 12'h1ee;
    rom[11922] = 12'h1ee;
    rom[11923] = 12'h1ee;
    rom[11924] = 12'h1ee;
    rom[11925] = 12'h1ee;
    rom[11926] = 12'h1ee;
    rom[11927] = 12'h1ee;
    rom[11928] = 12'h1ee;
    rom[11929] = 12'h000;
    rom[11930] = 12'h000;
    rom[11931] = 12'h000;
    rom[11932] = 12'h000;
    rom[11933] = 12'h000;
    rom[11934] = 12'h000;
    rom[11935] = 12'h000;
    rom[11936] = 12'h000;
    rom[11937] = 12'h000;
    rom[11938] = 12'h000;
    rom[11939] = 12'h000;
    rom[11940] = 12'h000;
    rom[11941] = 12'h000;
    rom[11942] = 12'h000;
    rom[11943] = 12'h000;
    rom[11944] = 12'h000;
    rom[11945] = 12'h000;
    rom[11946] = 12'h000;
    rom[11947] = 12'h000;
    rom[11948] = 12'h000;
    rom[11949] = 12'h000;
    rom[11950] = 12'h000;
    rom[11951] = 12'h000;
    rom[11952] = 12'h000;
    rom[11953] = 12'h000;
    rom[11954] = 12'h000;
    rom[11955] = 12'h000;
    rom[11956] = 12'h000;
    rom[11957] = 12'h000;
    rom[11958] = 12'h000;
    rom[11959] = 12'h000;
    rom[11960] = 12'h000;
    rom[11961] = 12'h000;
    rom[11962] = 12'h000;
    rom[11963] = 12'h000;
    rom[11964] = 12'h000;
    rom[11965] = 12'h000;
    rom[11966] = 12'h000;
    rom[11967] = 12'h000;
    rom[11968] = 12'h000;
    rom[11969] = 12'h000;
    rom[11970] = 12'h000;
    rom[11971] = 12'h000;
    rom[11972] = 12'h000;
    rom[11973] = 12'h000;
    rom[11974] = 12'h000;
    rom[11975] = 12'h000;
    rom[11976] = 12'h000;
    rom[11977] = 12'h000;
    rom[11978] = 12'h000;
    rom[11979] = 12'h000;
    rom[11980] = 12'h000;
    rom[11981] = 12'h000;
    rom[11982] = 12'h000;
    rom[11983] = 12'h000;
    rom[11984] = 12'h000;
    rom[11985] = 12'h000;
    rom[11986] = 12'h000;
    rom[11987] = 12'h000;
    rom[11988] = 12'h000;
    rom[11989] = 12'h000;
    rom[11990] = 12'h000;
    rom[11991] = 12'h000;
    rom[11992] = 12'h000;
    rom[11993] = 12'h000;
    rom[11994] = 12'h000;
    rom[11995] = 12'h000;
    rom[11996] = 12'h000;
    rom[11997] = 12'h000;
    rom[11998] = 12'h000;
    rom[11999] = 12'h000;
    rom[12000] = 12'h000;
    rom[12001] = 12'h000;
    rom[12002] = 12'h000;
    rom[12003] = 12'h000;
    rom[12004] = 12'h000;
    rom[12005] = 12'h000;
    rom[12006] = 12'h000;
    rom[12007] = 12'h3a2;
    rom[12008] = 12'h3a2;
    rom[12009] = 12'h3a2;
    rom[12010] = 12'h3a2;
    rom[12011] = 12'h3a2;
    rom[12012] = 12'h3a2;
    rom[12013] = 12'h3a2;
    rom[12014] = 12'h3a2;
    rom[12015] = 12'h3a2;
    rom[12016] = 12'h3a2;
    rom[12017] = 12'h3a2;
    rom[12018] = 12'h3a2;
    rom[12019] = 12'h3a2;
    rom[12020] = 12'h3a2;
    rom[12021] = 12'h3a2;
    rom[12022] = 12'h3a2;
    rom[12023] = 12'h3a2;
    rom[12024] = 12'h3a2;
    rom[12025] = 12'h000;
    rom[12026] = 12'h000;
    rom[12027] = 12'h000;
    rom[12028] = 12'h000;
    rom[12029] = 12'h000;
    rom[12030] = 12'h000;
    rom[12031] = 12'h000;
    rom[12032] = 12'h000;
    rom[12033] = 12'h000;
    rom[12034] = 12'h000;
    rom[12035] = 12'h000;
    rom[12036] = 12'h000;
    rom[12037] = 12'h000;
    rom[12038] = 12'h000;
    rom[12039] = 12'h000;
    rom[12040] = 12'h1ee;
    rom[12041] = 12'h1ee;
    rom[12042] = 12'h1ee;
    rom[12043] = 12'h1ee;
    rom[12044] = 12'h1ee;
    rom[12045] = 12'h1ee;
    rom[12046] = 12'h1ee;
    rom[12047] = 12'h1ee;
    rom[12048] = 12'h1ee;
    rom[12049] = 12'h1ee;
    rom[12050] = 12'h1ee;
    rom[12051] = 12'h1ee;
    rom[12052] = 12'h1ee;
    rom[12053] = 12'h1ee;
    rom[12054] = 12'h1ee;
    rom[12055] = 12'h1ee;
    rom[12056] = 12'h1ee;
    rom[12057] = 12'h1ee;
    rom[12058] = 12'h000;
    rom[12059] = 12'h000;
    rom[12060] = 12'h000;
    rom[12061] = 12'h000;
    rom[12062] = 12'h000;
    rom[12063] = 12'h000;
    rom[12064] = 12'h000;
    rom[12065] = 12'h000;
    rom[12066] = 12'h000;
    rom[12067] = 12'h000;
    rom[12068] = 12'h000;
    rom[12069] = 12'h000;
    rom[12070] = 12'h000;
    rom[12071] = 12'h000;
    rom[12072] = 12'h000;
    rom[12073] = 12'h000;
    rom[12074] = 12'h000;
    rom[12075] = 12'h000;
    rom[12076] = 12'h000;
    rom[12077] = 12'h000;
    rom[12078] = 12'h000;
    rom[12079] = 12'h000;
    rom[12080] = 12'h000;
    rom[12081] = 12'h000;
    rom[12082] = 12'h000;
    rom[12083] = 12'h000;
    rom[12084] = 12'h000;
    rom[12085] = 12'h000;
    rom[12086] = 12'h000;
    rom[12087] = 12'h000;
    rom[12088] = 12'h000;
    rom[12089] = 12'h000;
    rom[12090] = 12'h000;
    rom[12091] = 12'h000;
    rom[12092] = 12'h000;
    rom[12093] = 12'h000;
    rom[12094] = 12'h000;
    rom[12095] = 12'h000;
    rom[12096] = 12'h000;
    rom[12097] = 12'h000;
    rom[12098] = 12'h000;
    rom[12099] = 12'h000;
    rom[12100] = 12'h000;
    rom[12101] = 12'h000;
    rom[12102] = 12'h000;
    rom[12103] = 12'h000;
    rom[12104] = 12'h000;
    rom[12105] = 12'h000;
    rom[12106] = 12'h000;
    rom[12107] = 12'h000;
    rom[12108] = 12'h000;
    rom[12109] = 12'h000;
    rom[12110] = 12'h000;
    rom[12111] = 12'h000;
    rom[12112] = 12'h000;
    rom[12113] = 12'h000;
    rom[12114] = 12'h000;
    rom[12115] = 12'h000;
    rom[12116] = 12'h000;
    rom[12117] = 12'h000;
    rom[12118] = 12'h000;
    rom[12119] = 12'h000;
    rom[12120] = 12'h000;
    rom[12121] = 12'h000;
    rom[12122] = 12'h000;
    rom[12123] = 12'h000;
    rom[12124] = 12'h000;
    rom[12125] = 12'h000;
    rom[12126] = 12'h000;
    rom[12127] = 12'h000;
    rom[12128] = 12'h000;
    rom[12129] = 12'h000;
    rom[12130] = 12'h000;
    rom[12131] = 12'h000;
    rom[12132] = 12'h000;
    rom[12133] = 12'h000;
    rom[12134] = 12'h391;
    rom[12135] = 12'h3a2;
    rom[12136] = 12'h3a2;
    rom[12137] = 12'h3a2;
    rom[12138] = 12'h3a2;
    rom[12139] = 12'h3a2;
    rom[12140] = 12'h3a2;
    rom[12141] = 12'h3a2;
    rom[12142] = 12'h3a2;
    rom[12143] = 12'h3a2;
    rom[12144] = 12'h3a2;
    rom[12145] = 12'h3a2;
    rom[12146] = 12'h3a2;
    rom[12147] = 12'h3a2;
    rom[12148] = 12'h3a2;
    rom[12149] = 12'h3a2;
    rom[12150] = 12'h3a2;
    rom[12151] = 12'h3a2;
    rom[12152] = 12'h000;
    rom[12153] = 12'h000;
    rom[12154] = 12'h000;
    rom[12155] = 12'h000;
    rom[12156] = 12'h000;
    rom[12157] = 12'h000;
    rom[12158] = 12'h000;
    rom[12159] = 12'h000;
    rom[12160] = 12'h000;
    rom[12161] = 12'h000;
    rom[12162] = 12'h000;
    rom[12163] = 12'h000;
    rom[12164] = 12'h000;
    rom[12165] = 12'h000;
    rom[12166] = 12'h000;
    rom[12167] = 12'h000;
    rom[12168] = 12'h1ee;
    rom[12169] = 12'h1ee;
    rom[12170] = 12'h1ee;
    rom[12171] = 12'h1ee;
    rom[12172] = 12'h1ee;
    rom[12173] = 12'h1ee;
    rom[12174] = 12'h1ee;
    rom[12175] = 12'h1ee;
    rom[12176] = 12'h1ee;
    rom[12177] = 12'h1ee;
    rom[12178] = 12'h1ee;
    rom[12179] = 12'h1ee;
    rom[12180] = 12'h1ee;
    rom[12181] = 12'h1ee;
    rom[12182] = 12'h1ee;
    rom[12183] = 12'h1ee;
    rom[12184] = 12'h1ee;
    rom[12185] = 12'h1ee;
    rom[12186] = 12'h000;
    rom[12187] = 12'h000;
    rom[12188] = 12'h000;
    rom[12189] = 12'h000;
    rom[12190] = 12'h000;
    rom[12191] = 12'h000;
    rom[12192] = 12'h000;
    rom[12193] = 12'h000;
    rom[12194] = 12'h000;
    rom[12195] = 12'h000;
    rom[12196] = 12'h000;
    rom[12197] = 12'h000;
    rom[12198] = 12'h000;
    rom[12199] = 12'h000;
    rom[12200] = 12'h000;
    rom[12201] = 12'h000;
    rom[12202] = 12'h000;
    rom[12203] = 12'h000;
    rom[12204] = 12'h000;
    rom[12205] = 12'h000;
    rom[12206] = 12'h000;
    rom[12207] = 12'h000;
    rom[12208] = 12'h000;
    rom[12209] = 12'h000;
    rom[12210] = 12'h000;
    rom[12211] = 12'h000;
    rom[12212] = 12'h000;
    rom[12213] = 12'h000;
    rom[12214] = 12'h000;
    rom[12215] = 12'h000;
    rom[12216] = 12'h000;
    rom[12217] = 12'h000;
    rom[12218] = 12'h000;
    rom[12219] = 12'h000;
    rom[12220] = 12'h000;
    rom[12221] = 12'h000;
    rom[12222] = 12'h000;
    rom[12223] = 12'h000;
    rom[12224] = 12'h000;
    rom[12225] = 12'h000;
    rom[12226] = 12'h000;
    rom[12227] = 12'h000;
    rom[12228] = 12'h000;
    rom[12229] = 12'h000;
    rom[12230] = 12'h000;
    rom[12231] = 12'h000;
    rom[12232] = 12'h000;
    rom[12233] = 12'h000;
    rom[12234] = 12'h000;
    rom[12235] = 12'h000;
    rom[12236] = 12'h000;
    rom[12237] = 12'h000;
    rom[12238] = 12'h000;
    rom[12239] = 12'h000;
    rom[12240] = 12'h000;
    rom[12241] = 12'h000;
    rom[12242] = 12'h000;
    rom[12243] = 12'h000;
    rom[12244] = 12'h000;
    rom[12245] = 12'h000;
    rom[12246] = 12'h000;
    rom[12247] = 12'h000;
    rom[12248] = 12'h000;
    rom[12249] = 12'h000;
    rom[12250] = 12'h000;
    rom[12251] = 12'h000;
    rom[12252] = 12'h000;
    rom[12253] = 12'h000;
    rom[12254] = 12'h000;
    rom[12255] = 12'h000;
    rom[12256] = 12'h000;
    rom[12257] = 12'h000;
    rom[12258] = 12'h000;
    rom[12259] = 12'h000;
    rom[12260] = 12'h000;
    rom[12261] = 12'h000;
    rom[12262] = 12'h3a2;
    rom[12263] = 12'h3a2;
    rom[12264] = 12'h3a2;
    rom[12265] = 12'h3a2;
    rom[12266] = 12'h3a2;
    rom[12267] = 12'h3a2;
    rom[12268] = 12'h3a2;
    rom[12269] = 12'h3a2;
    rom[12270] = 12'h3a2;
    rom[12271] = 12'h3a2;
    rom[12272] = 12'h3a2;
    rom[12273] = 12'h3a2;
    rom[12274] = 12'h3a2;
    rom[12275] = 12'h3a2;
    rom[12276] = 12'h3a2;
    rom[12277] = 12'h3a2;
    rom[12278] = 12'h3a2;
    rom[12279] = 12'h3a2;
    rom[12280] = 12'h000;
    rom[12281] = 12'h000;
    rom[12282] = 12'h000;
    rom[12283] = 12'h000;
    rom[12284] = 12'h000;
    rom[12285] = 12'h000;
    rom[12286] = 12'h000;
    rom[12287] = 12'h000;
    rom[12288] = 12'h000;
    rom[12289] = 12'h000;
    rom[12290] = 12'h000;
    rom[12291] = 12'h000;
    rom[12292] = 12'h000;
    rom[12293] = 12'h000;
    rom[12294] = 12'h000;
    rom[12295] = 12'h000;
    rom[12296] = 12'h000;
    rom[12297] = 12'h1ee;
    rom[12298] = 12'h1ee;
    rom[12299] = 12'h1ee;
    rom[12300] = 12'h1ee;
    rom[12301] = 12'h1ee;
    rom[12302] = 12'h1ee;
    rom[12303] = 12'h1ee;
    rom[12304] = 12'h1ee;
    rom[12305] = 12'h1ee;
    rom[12306] = 12'h1ee;
    rom[12307] = 12'h1ee;
    rom[12308] = 12'h1ee;
    rom[12309] = 12'h1ee;
    rom[12310] = 12'h1ee;
    rom[12311] = 12'h1ef;
    rom[12312] = 12'h1ef;
    rom[12313] = 12'h1ef;
    rom[12314] = 12'h1ef;
    rom[12315] = 12'h000;
    rom[12316] = 12'h000;
    rom[12317] = 12'h000;
    rom[12318] = 12'h000;
    rom[12319] = 12'h000;
    rom[12320] = 12'h000;
    rom[12321] = 12'h000;
    rom[12322] = 12'h000;
    rom[12323] = 12'h000;
    rom[12324] = 12'h000;
    rom[12325] = 12'h000;
    rom[12326] = 12'h000;
    rom[12327] = 12'h000;
    rom[12328] = 12'h000;
    rom[12329] = 12'h000;
    rom[12330] = 12'h000;
    rom[12331] = 12'h000;
    rom[12332] = 12'h000;
    rom[12333] = 12'h000;
    rom[12334] = 12'h000;
    rom[12335] = 12'h000;
    rom[12336] = 12'h000;
    rom[12337] = 12'h000;
    rom[12338] = 12'h000;
    rom[12339] = 12'h000;
    rom[12340] = 12'h000;
    rom[12341] = 12'h000;
    rom[12342] = 12'h000;
    rom[12343] = 12'h000;
    rom[12344] = 12'h000;
    rom[12345] = 12'h000;
    rom[12346] = 12'h000;
    rom[12347] = 12'h000;
    rom[12348] = 12'h000;
    rom[12349] = 12'h000;
    rom[12350] = 12'h000;
    rom[12351] = 12'h000;
    rom[12352] = 12'h000;
    rom[12353] = 12'h000;
    rom[12354] = 12'h000;
    rom[12355] = 12'h000;
    rom[12356] = 12'h000;
    rom[12357] = 12'h000;
    rom[12358] = 12'h000;
    rom[12359] = 12'h000;
    rom[12360] = 12'h000;
    rom[12361] = 12'h000;
    rom[12362] = 12'h000;
    rom[12363] = 12'h000;
    rom[12364] = 12'h000;
    rom[12365] = 12'h000;
    rom[12366] = 12'h000;
    rom[12367] = 12'h000;
    rom[12368] = 12'h000;
    rom[12369] = 12'h000;
    rom[12370] = 12'h000;
    rom[12371] = 12'h000;
    rom[12372] = 12'h000;
    rom[12373] = 12'h000;
    rom[12374] = 12'h000;
    rom[12375] = 12'h000;
    rom[12376] = 12'h000;
    rom[12377] = 12'h000;
    rom[12378] = 12'h000;
    rom[12379] = 12'h000;
    rom[12380] = 12'h000;
    rom[12381] = 12'h000;
    rom[12382] = 12'h000;
    rom[12383] = 12'h000;
    rom[12384] = 12'h000;
    rom[12385] = 12'h000;
    rom[12386] = 12'h000;
    rom[12387] = 12'h000;
    rom[12388] = 12'h000;
    rom[12389] = 12'h3a2;
    rom[12390] = 12'h3a2;
    rom[12391] = 12'h3a2;
    rom[12392] = 12'h3a2;
    rom[12393] = 12'h3a2;
    rom[12394] = 12'h3a2;
    rom[12395] = 12'h3a2;
    rom[12396] = 12'h3a2;
    rom[12397] = 12'h3a2;
    rom[12398] = 12'h3a2;
    rom[12399] = 12'h3a2;
    rom[12400] = 12'h3a2;
    rom[12401] = 12'h3a2;
    rom[12402] = 12'h3a2;
    rom[12403] = 12'h3a2;
    rom[12404] = 12'h3a2;
    rom[12405] = 12'h3a2;
    rom[12406] = 12'h3a2;
    rom[12407] = 12'h000;
    rom[12408] = 12'h000;
    rom[12409] = 12'h000;
    rom[12410] = 12'h000;
    rom[12411] = 12'h000;
    rom[12412] = 12'h000;
    rom[12413] = 12'h000;
    rom[12414] = 12'h000;
    rom[12415] = 12'h000;
    rom[12416] = 12'h000;
    rom[12417] = 12'h000;
    rom[12418] = 12'h000;
    rom[12419] = 12'h000;
    rom[12420] = 12'h000;
    rom[12421] = 12'h000;
    rom[12422] = 12'h000;
    rom[12423] = 12'h000;
    rom[12424] = 12'h000;
    rom[12425] = 12'h1dd;
    rom[12426] = 12'h1ee;
    rom[12427] = 12'h1ee;
    rom[12428] = 12'h1ee;
    rom[12429] = 12'h1ee;
    rom[12430] = 12'h1ee;
    rom[12431] = 12'h1ee;
    rom[12432] = 12'h1ee;
    rom[12433] = 12'h1ee;
    rom[12434] = 12'h1ee;
    rom[12435] = 12'h1ee;
    rom[12436] = 12'h1ef;
    rom[12437] = 12'h1ef;
    rom[12438] = 12'h1ef;
    rom[12439] = 12'h1ef;
    rom[12440] = 12'h1ef;
    rom[12441] = 12'h1ef;
    rom[12442] = 12'h1ef;
    rom[12443] = 12'h1ef;
    rom[12444] = 12'h000;
    rom[12445] = 12'h000;
    rom[12446] = 12'h000;
    rom[12447] = 12'h000;
    rom[12448] = 12'h000;
    rom[12449] = 12'h000;
    rom[12450] = 12'h000;
    rom[12451] = 12'h000;
    rom[12452] = 12'h000;
    rom[12453] = 12'h000;
    rom[12454] = 12'h000;
    rom[12455] = 12'h000;
    rom[12456] = 12'h000;
    rom[12457] = 12'h000;
    rom[12458] = 12'h000;
    rom[12459] = 12'h000;
    rom[12460] = 12'h000;
    rom[12461] = 12'h000;
    rom[12462] = 12'h000;
    rom[12463] = 12'h000;
    rom[12464] = 12'h000;
    rom[12465] = 12'h000;
    rom[12466] = 12'h000;
    rom[12467] = 12'h000;
    rom[12468] = 12'h000;
    rom[12469] = 12'h000;
    rom[12470] = 12'h000;
    rom[12471] = 12'h000;
    rom[12472] = 12'h000;
    rom[12473] = 12'h000;
    rom[12474] = 12'h000;
    rom[12475] = 12'h000;
    rom[12476] = 12'h000;
    rom[12477] = 12'h000;
    rom[12478] = 12'h000;
    rom[12479] = 12'h000;
    rom[12480] = 12'h000;
    rom[12481] = 12'h000;
    rom[12482] = 12'h000;
    rom[12483] = 12'h000;
    rom[12484] = 12'h000;
    rom[12485] = 12'h000;
    rom[12486] = 12'h000;
    rom[12487] = 12'h000;
    rom[12488] = 12'h000;
    rom[12489] = 12'h000;
    rom[12490] = 12'h000;
    rom[12491] = 12'h000;
    rom[12492] = 12'h000;
    rom[12493] = 12'h000;
    rom[12494] = 12'h000;
    rom[12495] = 12'h000;
    rom[12496] = 12'h000;
    rom[12497] = 12'h000;
    rom[12498] = 12'h000;
    rom[12499] = 12'h000;
    rom[12500] = 12'h000;
    rom[12501] = 12'h000;
    rom[12502] = 12'h000;
    rom[12503] = 12'h000;
    rom[12504] = 12'h000;
    rom[12505] = 12'h000;
    rom[12506] = 12'h000;
    rom[12507] = 12'h000;
    rom[12508] = 12'h000;
    rom[12509] = 12'h000;
    rom[12510] = 12'h000;
    rom[12511] = 12'h000;
    rom[12512] = 12'h000;
    rom[12513] = 12'h000;
    rom[12514] = 12'h000;
    rom[12515] = 12'h000;
    rom[12516] = 12'h3a2;
    rom[12517] = 12'h3a2;
    rom[12518] = 12'h3a2;
    rom[12519] = 12'h3a2;
    rom[12520] = 12'h3a2;
    rom[12521] = 12'h3a2;
    rom[12522] = 12'h3a2;
    rom[12523] = 12'h3a2;
    rom[12524] = 12'h3a2;
    rom[12525] = 12'h3a2;
    rom[12526] = 12'h3a2;
    rom[12527] = 12'h3a2;
    rom[12528] = 12'h3a2;
    rom[12529] = 12'h3a2;
    rom[12530] = 12'h3a2;
    rom[12531] = 12'h3a2;
    rom[12532] = 12'h3a2;
    rom[12533] = 12'h3a2;
    rom[12534] = 12'h3a2;
    rom[12535] = 12'h000;
    rom[12536] = 12'h000;
    rom[12537] = 12'h000;
    rom[12538] = 12'h000;
    rom[12539] = 12'h000;
    rom[12540] = 12'h000;
    rom[12541] = 12'h000;
    rom[12542] = 12'h000;
    rom[12543] = 12'h000;
    rom[12544] = 12'h000;
    rom[12545] = 12'h000;
    rom[12546] = 12'h000;
    rom[12547] = 12'h000;
    rom[12548] = 12'h000;
    rom[12549] = 12'h000;
    rom[12550] = 12'h000;
    rom[12551] = 12'h000;
    rom[12552] = 12'h000;
    rom[12553] = 12'h000;
    rom[12554] = 12'h1ee;
    rom[12555] = 12'h1ee;
    rom[12556] = 12'h1ee;
    rom[12557] = 12'h1ee;
    rom[12558] = 12'h1ee;
    rom[12559] = 12'h1ee;
    rom[12560] = 12'h1ee;
    rom[12561] = 12'h1ee;
    rom[12562] = 12'h1ef;
    rom[12563] = 12'h1ef;
    rom[12564] = 12'h1ef;
    rom[12565] = 12'h1ef;
    rom[12566] = 12'h1ef;
    rom[12567] = 12'h1ef;
    rom[12568] = 12'h1ef;
    rom[12569] = 12'h1ef;
    rom[12570] = 12'h1ef;
    rom[12571] = 12'h1ef;
    rom[12572] = 12'h1ef;
    rom[12573] = 12'h000;
    rom[12574] = 12'h000;
    rom[12575] = 12'h000;
    rom[12576] = 12'h000;
    rom[12577] = 12'h000;
    rom[12578] = 12'h000;
    rom[12579] = 12'h000;
    rom[12580] = 12'h000;
    rom[12581] = 12'h000;
    rom[12582] = 12'h000;
    rom[12583] = 12'h000;
    rom[12584] = 12'h000;
    rom[12585] = 12'h000;
    rom[12586] = 12'h000;
    rom[12587] = 12'h000;
    rom[12588] = 12'h000;
    rom[12589] = 12'h000;
    rom[12590] = 12'h000;
    rom[12591] = 12'h000;
    rom[12592] = 12'h000;
    rom[12593] = 12'h000;
    rom[12594] = 12'h000;
    rom[12595] = 12'h000;
    rom[12596] = 12'h000;
    rom[12597] = 12'h000;
    rom[12598] = 12'h000;
    rom[12599] = 12'h000;
    rom[12600] = 12'h000;
    rom[12601] = 12'h000;
    rom[12602] = 12'h000;
    rom[12603] = 12'h000;
    rom[12604] = 12'h000;
    rom[12605] = 12'h000;
    rom[12606] = 12'h000;
    rom[12607] = 12'h000;
    rom[12608] = 12'h000;
    rom[12609] = 12'h000;
    rom[12610] = 12'h000;
    rom[12611] = 12'h000;
    rom[12612] = 12'h000;
    rom[12613] = 12'h000;
    rom[12614] = 12'h000;
    rom[12615] = 12'h000;
    rom[12616] = 12'h000;
    rom[12617] = 12'h000;
    rom[12618] = 12'h000;
    rom[12619] = 12'h000;
    rom[12620] = 12'h000;
    rom[12621] = 12'h000;
    rom[12622] = 12'h000;
    rom[12623] = 12'h000;
    rom[12624] = 12'h000;
    rom[12625] = 12'h000;
    rom[12626] = 12'h000;
    rom[12627] = 12'h000;
    rom[12628] = 12'h000;
    rom[12629] = 12'h000;
    rom[12630] = 12'h000;
    rom[12631] = 12'h000;
    rom[12632] = 12'h000;
    rom[12633] = 12'h000;
    rom[12634] = 12'h000;
    rom[12635] = 12'h000;
    rom[12636] = 12'h000;
    rom[12637] = 12'h000;
    rom[12638] = 12'h000;
    rom[12639] = 12'h000;
    rom[12640] = 12'h000;
    rom[12641] = 12'h000;
    rom[12642] = 12'h000;
    rom[12643] = 12'h3a2;
    rom[12644] = 12'h3a2;
    rom[12645] = 12'h3a2;
    rom[12646] = 12'h3a2;
    rom[12647] = 12'h3a2;
    rom[12648] = 12'h3a2;
    rom[12649] = 12'h3a2;
    rom[12650] = 12'h3a2;
    rom[12651] = 12'h3a2;
    rom[12652] = 12'h3a2;
    rom[12653] = 12'h3a2;
    rom[12654] = 12'h3a2;
    rom[12655] = 12'h3a2;
    rom[12656] = 12'h3a2;
    rom[12657] = 12'h3a2;
    rom[12658] = 12'h3a2;
    rom[12659] = 12'h3a2;
    rom[12660] = 12'h3a2;
    rom[12661] = 12'h3a2;
    rom[12662] = 12'h000;
    rom[12663] = 12'h000;
    rom[12664] = 12'h000;
    rom[12665] = 12'h000;
    rom[12666] = 12'h000;
    rom[12667] = 12'h000;
    rom[12668] = 12'h000;
    rom[12669] = 12'h000;
    rom[12670] = 12'h000;
    rom[12671] = 12'h000;
    rom[12672] = 12'h000;
    rom[12673] = 12'h000;
    rom[12674] = 12'h000;
    rom[12675] = 12'h000;
    rom[12676] = 12'h000;
    rom[12677] = 12'h000;
    rom[12678] = 12'h000;
    rom[12679] = 12'h000;
    rom[12680] = 12'h000;
    rom[12681] = 12'h000;
    rom[12682] = 12'h000;
    rom[12683] = 12'h1ee;
    rom[12684] = 12'h1ee;
    rom[12685] = 12'h1ee;
    rom[12686] = 12'h1ee;
    rom[12687] = 12'h1ef;
    rom[12688] = 12'h1ef;
    rom[12689] = 12'h1ef;
    rom[12690] = 12'h1ef;
    rom[12691] = 12'h1ef;
    rom[12692] = 12'h1ef;
    rom[12693] = 12'h1ef;
    rom[12694] = 12'h1ef;
    rom[12695] = 12'h1ef;
    rom[12696] = 12'h1ef;
    rom[12697] = 12'h1ef;
    rom[12698] = 12'h1ef;
    rom[12699] = 12'h1ef;
    rom[12700] = 12'h1ef;
    rom[12701] = 12'h1ef;
    rom[12702] = 12'h000;
    rom[12703] = 12'h000;
    rom[12704] = 12'h000;
    rom[12705] = 12'h000;
    rom[12706] = 12'h000;
    rom[12707] = 12'h000;
    rom[12708] = 12'h000;
    rom[12709] = 12'h000;
    rom[12710] = 12'h000;
    rom[12711] = 12'h000;
    rom[12712] = 12'h000;
    rom[12713] = 12'h000;
    rom[12714] = 12'h000;
    rom[12715] = 12'h000;
    rom[12716] = 12'h000;
    rom[12717] = 12'h000;
    rom[12718] = 12'h000;
    rom[12719] = 12'h000;
    rom[12720] = 12'h000;
    rom[12721] = 12'h000;
    rom[12722] = 12'h000;
    rom[12723] = 12'h000;
    rom[12724] = 12'h000;
    rom[12725] = 12'h000;
    rom[12726] = 12'h000;
    rom[12727] = 12'h000;
    rom[12728] = 12'h000;
    rom[12729] = 12'h000;
    rom[12730] = 12'h000;
    rom[12731] = 12'h000;
    rom[12732] = 12'h000;
    rom[12733] = 12'h000;
    rom[12734] = 12'h000;
    rom[12735] = 12'h000;
    rom[12736] = 12'h000;
    rom[12737] = 12'h000;
    rom[12738] = 12'h000;
    rom[12739] = 12'h000;
    rom[12740] = 12'h000;
    rom[12741] = 12'h000;
    rom[12742] = 12'h000;
    rom[12743] = 12'h000;
    rom[12744] = 12'h000;
    rom[12745] = 12'h000;
    rom[12746] = 12'h000;
    rom[12747] = 12'h000;
    rom[12748] = 12'h000;
    rom[12749] = 12'h000;
    rom[12750] = 12'h000;
    rom[12751] = 12'h000;
    rom[12752] = 12'h000;
    rom[12753] = 12'h000;
    rom[12754] = 12'h000;
    rom[12755] = 12'h000;
    rom[12756] = 12'h000;
    rom[12757] = 12'h000;
    rom[12758] = 12'h000;
    rom[12759] = 12'h000;
    rom[12760] = 12'h000;
    rom[12761] = 12'h000;
    rom[12762] = 12'h000;
    rom[12763] = 12'h000;
    rom[12764] = 12'h000;
    rom[12765] = 12'h000;
    rom[12766] = 12'h000;
    rom[12767] = 12'h000;
    rom[12768] = 12'h000;
    rom[12769] = 12'h000;
    rom[12770] = 12'h3a2;
    rom[12771] = 12'h3a2;
    rom[12772] = 12'h3a2;
    rom[12773] = 12'h3a2;
    rom[12774] = 12'h3a2;
    rom[12775] = 12'h3a2;
    rom[12776] = 12'h3a2;
    rom[12777] = 12'h3a2;
    rom[12778] = 12'h3a2;
    rom[12779] = 12'h3a2;
    rom[12780] = 12'h3a2;
    rom[12781] = 12'h3a2;
    rom[12782] = 12'h3a2;
    rom[12783] = 12'h3a2;
    rom[12784] = 12'h3a2;
    rom[12785] = 12'h3a2;
    rom[12786] = 12'h3a2;
    rom[12787] = 12'h3a2;
    rom[12788] = 12'h3a2;
    rom[12789] = 12'h000;
    rom[12790] = 12'h000;
    rom[12791] = 12'h000;
    rom[12792] = 12'h000;
    rom[12793] = 12'h000;
    rom[12794] = 12'h000;
    rom[12795] = 12'h000;
    rom[12796] = 12'h000;
    rom[12797] = 12'h000;
    rom[12798] = 12'h000;
    rom[12799] = 12'h000;
    rom[12800] = 12'h000;
    rom[12801] = 12'h000;
    rom[12802] = 12'h000;
    rom[12803] = 12'h000;
    rom[12804] = 12'h000;
    rom[12805] = 12'h000;
    rom[12806] = 12'h000;
    rom[12807] = 12'h000;
    rom[12808] = 12'h000;
    rom[12809] = 12'h000;
    rom[12810] = 12'h000;
    rom[12811] = 12'h1ee;
    rom[12812] = 12'h1ef;
    rom[12813] = 12'h1ef;
    rom[12814] = 12'h1ef;
    rom[12815] = 12'h1ef;
    rom[12816] = 12'h1ef;
    rom[12817] = 12'h1ef;
    rom[12818] = 12'h1ef;
    rom[12819] = 12'h1ef;
    rom[12820] = 12'h1ef;
    rom[12821] = 12'h1ef;
    rom[12822] = 12'h1ef;
    rom[12823] = 12'h1ef;
    rom[12824] = 12'h1ef;
    rom[12825] = 12'h1ef;
    rom[12826] = 12'h1ef;
    rom[12827] = 12'h1ef;
    rom[12828] = 12'h1ef;
    rom[12829] = 12'h1ef;
    rom[12830] = 12'h1ef;
    rom[12831] = 12'h000;
    rom[12832] = 12'h000;
    rom[12833] = 12'h000;
    rom[12834] = 12'h000;
    rom[12835] = 12'h000;
    rom[12836] = 12'h000;
    rom[12837] = 12'h000;
    rom[12838] = 12'h000;
    rom[12839] = 12'h000;
    rom[12840] = 12'h000;
    rom[12841] = 12'h000;
    rom[12842] = 12'h000;
    rom[12843] = 12'h000;
    rom[12844] = 12'h000;
    rom[12845] = 12'h000;
    rom[12846] = 12'h000;
    rom[12847] = 12'h000;
    rom[12848] = 12'h000;
    rom[12849] = 12'h000;
    rom[12850] = 12'h000;
    rom[12851] = 12'h000;
    rom[12852] = 12'h000;
    rom[12853] = 12'h000;
    rom[12854] = 12'h000;
    rom[12855] = 12'h000;
    rom[12856] = 12'h000;
    rom[12857] = 12'h000;
    rom[12858] = 12'h000;
    rom[12859] = 12'h000;
    rom[12860] = 12'h000;
    rom[12861] = 12'h000;
    rom[12862] = 12'h000;
    rom[12863] = 12'h000;
    rom[12864] = 12'h000;
    rom[12865] = 12'h000;
    rom[12866] = 12'h000;
    rom[12867] = 12'h000;
    rom[12868] = 12'h000;
    rom[12869] = 12'h000;
    rom[12870] = 12'h000;
    rom[12871] = 12'h000;
    rom[12872] = 12'h000;
    rom[12873] = 12'h000;
    rom[12874] = 12'h000;
    rom[12875] = 12'h000;
    rom[12876] = 12'h000;
    rom[12877] = 12'h000;
    rom[12878] = 12'h000;
    rom[12879] = 12'h000;
    rom[12880] = 12'h000;
    rom[12881] = 12'h000;
    rom[12882] = 12'h000;
    rom[12883] = 12'h000;
    rom[12884] = 12'h000;
    rom[12885] = 12'h000;
    rom[12886] = 12'h000;
    rom[12887] = 12'h000;
    rom[12888] = 12'h000;
    rom[12889] = 12'h000;
    rom[12890] = 12'h000;
    rom[12891] = 12'h000;
    rom[12892] = 12'h000;
    rom[12893] = 12'h000;
    rom[12894] = 12'h000;
    rom[12895] = 12'h000;
    rom[12896] = 12'h000;
    rom[12897] = 12'h3a2;
    rom[12898] = 12'h3a2;
    rom[12899] = 12'h3a2;
    rom[12900] = 12'h3a2;
    rom[12901] = 12'h3a2;
    rom[12902] = 12'h3a2;
    rom[12903] = 12'h3a2;
    rom[12904] = 12'h3a2;
    rom[12905] = 12'h3a2;
    rom[12906] = 12'h3a2;
    rom[12907] = 12'h3a2;
    rom[12908] = 12'h3a2;
    rom[12909] = 12'h3a2;
    rom[12910] = 12'h3a2;
    rom[12911] = 12'h3a2;
    rom[12912] = 12'h3a2;
    rom[12913] = 12'h3a2;
    rom[12914] = 12'h3a2;
    rom[12915] = 12'h3a2;
    rom[12916] = 12'h3a2;
    rom[12917] = 12'h000;
    rom[12918] = 12'h000;
    rom[12919] = 12'h000;
    rom[12920] = 12'h000;
    rom[12921] = 12'h000;
    rom[12922] = 12'h000;
    rom[12923] = 12'h000;
    rom[12924] = 12'h000;
    rom[12925] = 12'h000;
    rom[12926] = 12'h000;
    rom[12927] = 12'h000;
    rom[12928] = 12'h000;
    rom[12929] = 12'h000;
    rom[12930] = 12'h000;
    rom[12931] = 12'h000;
    rom[12932] = 12'h000;
    rom[12933] = 12'h000;
    rom[12934] = 12'h000;
    rom[12935] = 12'h000;
    rom[12936] = 12'h000;
    rom[12937] = 12'h000;
    rom[12938] = 12'h000;
    rom[12939] = 12'h000;
    rom[12940] = 12'h1ef;
    rom[12941] = 12'h1ef;
    rom[12942] = 12'h1ef;
    rom[12943] = 12'h1ef;
    rom[12944] = 12'h1ef;
    rom[12945] = 12'h1ef;
    rom[12946] = 12'h1ef;
    rom[12947] = 12'h1ef;
    rom[12948] = 12'h1ef;
    rom[12949] = 12'h1ef;
    rom[12950] = 12'h1ef;
    rom[12951] = 12'h1ef;
    rom[12952] = 12'h1ef;
    rom[12953] = 12'h1ef;
    rom[12954] = 12'h1ef;
    rom[12955] = 12'h1ef;
    rom[12956] = 12'h1ef;
    rom[12957] = 12'h1ef;
    rom[12958] = 12'h1ef;
    rom[12959] = 12'h1ef;
    rom[12960] = 12'h000;
    rom[12961] = 12'h000;
    rom[12962] = 12'h000;
    rom[12963] = 12'h000;
    rom[12964] = 12'h000;
    rom[12965] = 12'h000;
    rom[12966] = 12'h000;
    rom[12967] = 12'h000;
    rom[12968] = 12'h000;
    rom[12969] = 12'h000;
    rom[12970] = 12'h000;
    rom[12971] = 12'h000;
    rom[12972] = 12'h000;
    rom[12973] = 12'h000;
    rom[12974] = 12'h000;
    rom[12975] = 12'h000;
    rom[12976] = 12'h000;
    rom[12977] = 12'h000;
    rom[12978] = 12'h000;
    rom[12979] = 12'h000;
    rom[12980] = 12'h000;
    rom[12981] = 12'h000;
    rom[12982] = 12'h000;
    rom[12983] = 12'h000;
    rom[12984] = 12'h000;
    rom[12985] = 12'h000;
    rom[12986] = 12'h000;
    rom[12987] = 12'h000;
    rom[12988] = 12'h000;
    rom[12989] = 12'h000;
    rom[12990] = 12'h000;
    rom[12991] = 12'h000;
    rom[12992] = 12'h000;
    rom[12993] = 12'h000;
    rom[12994] = 12'h000;
    rom[12995] = 12'h000;
    rom[12996] = 12'h000;
    rom[12997] = 12'h000;
    rom[12998] = 12'h000;
    rom[12999] = 12'h000;
    rom[13000] = 12'h000;
    rom[13001] = 12'h000;
    rom[13002] = 12'h000;
    rom[13003] = 12'h000;
    rom[13004] = 12'h000;
    rom[13005] = 12'h000;
    rom[13006] = 12'h000;
    rom[13007] = 12'h000;
    rom[13008] = 12'h000;
    rom[13009] = 12'h000;
    rom[13010] = 12'h000;
    rom[13011] = 12'h000;
    rom[13012] = 12'h000;
    rom[13013] = 12'h000;
    rom[13014] = 12'h000;
    rom[13015] = 12'h000;
    rom[13016] = 12'h000;
    rom[13017] = 12'h000;
    rom[13018] = 12'h000;
    rom[13019] = 12'h000;
    rom[13020] = 12'h000;
    rom[13021] = 12'h000;
    rom[13022] = 12'h000;
    rom[13023] = 12'h3a2;
    rom[13024] = 12'h3a2;
    rom[13025] = 12'h3a2;
    rom[13026] = 12'h3a2;
    rom[13027] = 12'h3a2;
    rom[13028] = 12'h3a2;
    rom[13029] = 12'h3a2;
    rom[13030] = 12'h3a2;
    rom[13031] = 12'h3a2;
    rom[13032] = 12'h3a2;
    rom[13033] = 12'h3a2;
    rom[13034] = 12'h3a2;
    rom[13035] = 12'h3a2;
    rom[13036] = 12'h3a2;
    rom[13037] = 12'h3a2;
    rom[13038] = 12'h3a2;
    rom[13039] = 12'h3a2;
    rom[13040] = 12'h3a2;
    rom[13041] = 12'h3a2;
    rom[13042] = 12'h3a2;
    rom[13043] = 12'h3a2;
    rom[13044] = 12'h000;
    rom[13045] = 12'h000;
    rom[13046] = 12'h000;
    rom[13047] = 12'h000;
    rom[13048] = 12'h000;
    rom[13049] = 12'h000;
    rom[13050] = 12'h000;
    rom[13051] = 12'h000;
    rom[13052] = 12'h000;
    rom[13053] = 12'h000;
    rom[13054] = 12'h000;
    rom[13055] = 12'h000;
    rom[13056] = 12'h000;
    rom[13057] = 12'h000;
    rom[13058] = 12'h000;
    rom[13059] = 12'h000;
    rom[13060] = 12'h000;
    rom[13061] = 12'h000;
    rom[13062] = 12'h000;
    rom[13063] = 12'h000;
    rom[13064] = 12'h000;
    rom[13065] = 12'h000;
    rom[13066] = 12'h000;
    rom[13067] = 12'h000;
    rom[13068] = 12'h000;
    rom[13069] = 12'h1ef;
    rom[13070] = 12'h1ef;
    rom[13071] = 12'h1ef;
    rom[13072] = 12'h1ef;
    rom[13073] = 12'h1ef;
    rom[13074] = 12'h1ef;
    rom[13075] = 12'h1ef;
    rom[13076] = 12'h1ef;
    rom[13077] = 12'h1ef;
    rom[13078] = 12'h1ef;
    rom[13079] = 12'h1ef;
    rom[13080] = 12'h1ef;
    rom[13081] = 12'h1ef;
    rom[13082] = 12'h1ef;
    rom[13083] = 12'h1ef;
    rom[13084] = 12'h1ef;
    rom[13085] = 12'h1ef;
    rom[13086] = 12'h1ef;
    rom[13087] = 12'h1ef;
    rom[13088] = 12'h1ee;
    rom[13089] = 12'h1ee;
    rom[13090] = 12'h000;
    rom[13091] = 12'h000;
    rom[13092] = 12'h000;
    rom[13093] = 12'h000;
    rom[13094] = 12'h000;
    rom[13095] = 12'h000;
    rom[13096] = 12'h000;
    rom[13097] = 12'h000;
    rom[13098] = 12'h000;
    rom[13099] = 12'h000;
    rom[13100] = 12'h000;
    rom[13101] = 12'h000;
    rom[13102] = 12'h000;
    rom[13103] = 12'h000;
    rom[13104] = 12'h000;
    rom[13105] = 12'h000;
    rom[13106] = 12'h000;
    rom[13107] = 12'h000;
    rom[13108] = 12'h000;
    rom[13109] = 12'h000;
    rom[13110] = 12'h000;
    rom[13111] = 12'h000;
    rom[13112] = 12'h000;
    rom[13113] = 12'h000;
    rom[13114] = 12'h000;
    rom[13115] = 12'h000;
    rom[13116] = 12'h000;
    rom[13117] = 12'h000;
    rom[13118] = 12'h000;
    rom[13119] = 12'h000;
    rom[13120] = 12'h000;
    rom[13121] = 12'h000;
    rom[13122] = 12'h000;
    rom[13123] = 12'h000;
    rom[13124] = 12'h000;
    rom[13125] = 12'h000;
    rom[13126] = 12'h000;
    rom[13127] = 12'h000;
    rom[13128] = 12'h000;
    rom[13129] = 12'h000;
    rom[13130] = 12'h000;
    rom[13131] = 12'h000;
    rom[13132] = 12'h000;
    rom[13133] = 12'h000;
    rom[13134] = 12'h000;
    rom[13135] = 12'h000;
    rom[13136] = 12'h000;
    rom[13137] = 12'h000;
    rom[13138] = 12'h000;
    rom[13139] = 12'h000;
    rom[13140] = 12'h000;
    rom[13141] = 12'h000;
    rom[13142] = 12'h000;
    rom[13143] = 12'h000;
    rom[13144] = 12'h000;
    rom[13145] = 12'h000;
    rom[13146] = 12'h000;
    rom[13147] = 12'h000;
    rom[13148] = 12'h000;
    rom[13149] = 12'h000;
    rom[13150] = 12'h3a3;
    rom[13151] = 12'h3a2;
    rom[13152] = 12'h3a2;
    rom[13153] = 12'h3a2;
    rom[13154] = 12'h3a2;
    rom[13155] = 12'h3a2;
    rom[13156] = 12'h3a2;
    rom[13157] = 12'h3a2;
    rom[13158] = 12'h3a2;
    rom[13159] = 12'h3a2;
    rom[13160] = 12'h3a2;
    rom[13161] = 12'h3a2;
    rom[13162] = 12'h3a2;
    rom[13163] = 12'h3a2;
    rom[13164] = 12'h3a2;
    rom[13165] = 12'h3a2;
    rom[13166] = 12'h3a2;
    rom[13167] = 12'h3a2;
    rom[13168] = 12'h3a2;
    rom[13169] = 12'h3a2;
    rom[13170] = 12'h3a2;
    rom[13171] = 12'h000;
    rom[13172] = 12'h000;
    rom[13173] = 12'h000;
    rom[13174] = 12'h000;
    rom[13175] = 12'h000;
    rom[13176] = 12'h000;
    rom[13177] = 12'h000;
    rom[13178] = 12'h000;
    rom[13179] = 12'h000;
    rom[13180] = 12'h000;
    rom[13181] = 12'h000;
    rom[13182] = 12'h000;
    rom[13183] = 12'h000;
    rom[13184] = 12'h000;
    rom[13185] = 12'h000;
    rom[13186] = 12'h000;
    rom[13187] = 12'h000;
    rom[13188] = 12'h000;
    rom[13189] = 12'h000;
    rom[13190] = 12'h000;
    rom[13191] = 12'h000;
    rom[13192] = 12'h000;
    rom[13193] = 12'h000;
    rom[13194] = 12'h000;
    rom[13195] = 12'h000;
    rom[13196] = 12'h000;
    rom[13197] = 12'h000;
    rom[13198] = 12'h1ef;
    rom[13199] = 12'h1ef;
    rom[13200] = 12'h1ef;
    rom[13201] = 12'h1ef;
    rom[13202] = 12'h1ef;
    rom[13203] = 12'h1ef;
    rom[13204] = 12'h1ef;
    rom[13205] = 12'h1ef;
    rom[13206] = 12'h1ef;
    rom[13207] = 12'h1ef;
    rom[13208] = 12'h1ef;
    rom[13209] = 12'h1ef;
    rom[13210] = 12'h1ef;
    rom[13211] = 12'h1ef;
    rom[13212] = 12'h1ef;
    rom[13213] = 12'h1ef;
    rom[13214] = 12'h1ef;
    rom[13215] = 12'h1ee;
    rom[13216] = 12'h1ee;
    rom[13217] = 12'h1ee;
    rom[13218] = 12'h1ee;
    rom[13219] = 12'h000;
    rom[13220] = 12'h000;
    rom[13221] = 12'h000;
    rom[13222] = 12'h000;
    rom[13223] = 12'h000;
    rom[13224] = 12'h000;
    rom[13225] = 12'h000;
    rom[13226] = 12'h000;
    rom[13227] = 12'h000;
    rom[13228] = 12'h000;
    rom[13229] = 12'h000;
    rom[13230] = 12'h000;
    rom[13231] = 12'h000;
    rom[13232] = 12'h000;
    rom[13233] = 12'h000;
    rom[13234] = 12'h000;
    rom[13235] = 12'h000;
    rom[13236] = 12'h000;
    rom[13237] = 12'h000;
    rom[13238] = 12'h000;
    rom[13239] = 12'h000;
    rom[13240] = 12'h000;
    rom[13241] = 12'h000;
    rom[13242] = 12'h000;
    rom[13243] = 12'h000;
    rom[13244] = 12'h000;
    rom[13245] = 12'h000;
    rom[13246] = 12'h000;
    rom[13247] = 12'h000;
    rom[13248] = 12'h000;
    rom[13249] = 12'h000;
    rom[13250] = 12'h000;
    rom[13251] = 12'h000;
    rom[13252] = 12'h000;
    rom[13253] = 12'h000;
    rom[13254] = 12'h000;
    rom[13255] = 12'h000;
    rom[13256] = 12'h000;
    rom[13257] = 12'h000;
    rom[13258] = 12'h000;
    rom[13259] = 12'h000;
    rom[13260] = 12'h000;
    rom[13261] = 12'h000;
    rom[13262] = 12'h000;
    rom[13263] = 12'h000;
    rom[13264] = 12'h000;
    rom[13265] = 12'h000;
    rom[13266] = 12'h000;
    rom[13267] = 12'h000;
    rom[13268] = 12'h000;
    rom[13269] = 12'h000;
    rom[13270] = 12'h000;
    rom[13271] = 12'h000;
    rom[13272] = 12'h000;
    rom[13273] = 12'h000;
    rom[13274] = 12'h000;
    rom[13275] = 12'h000;
    rom[13276] = 12'h000;
    rom[13277] = 12'h3a3;
    rom[13278] = 12'h3a3;
    rom[13279] = 12'h3a2;
    rom[13280] = 12'h3a2;
    rom[13281] = 12'h3a2;
    rom[13282] = 12'h3a2;
    rom[13283] = 12'h3a2;
    rom[13284] = 12'h3a2;
    rom[13285] = 12'h3a2;
    rom[13286] = 12'h3a2;
    rom[13287] = 12'h3a2;
    rom[13288] = 12'h3a2;
    rom[13289] = 12'h3a2;
    rom[13290] = 12'h3a2;
    rom[13291] = 12'h3a2;
    rom[13292] = 12'h3a2;
    rom[13293] = 12'h3a2;
    rom[13294] = 12'h3a2;
    rom[13295] = 12'h3a2;
    rom[13296] = 12'h3a2;
    rom[13297] = 12'h3a2;
    rom[13298] = 12'h0f0;
    rom[13299] = 12'h000;
    rom[13300] = 12'h000;
    rom[13301] = 12'h000;
    rom[13302] = 12'h000;
    rom[13303] = 12'h000;
    rom[13304] = 12'h000;
    rom[13305] = 12'h000;
    rom[13306] = 12'h000;
    rom[13307] = 12'h000;
    rom[13308] = 12'h000;
    rom[13309] = 12'h000;
    rom[13310] = 12'h000;
    rom[13311] = 12'h000;
    rom[13312] = 12'h000;
    rom[13313] = 12'h000;
    rom[13314] = 12'h000;
    rom[13315] = 12'h000;
    rom[13316] = 12'h000;
    rom[13317] = 12'h000;
    rom[13318] = 12'h000;
    rom[13319] = 12'h000;
    rom[13320] = 12'h000;
    rom[13321] = 12'h000;
    rom[13322] = 12'h000;
    rom[13323] = 12'h000;
    rom[13324] = 12'h000;
    rom[13325] = 12'h000;
    rom[13326] = 12'h1de;
    rom[13327] = 12'h1ef;
    rom[13328] = 12'h1ef;
    rom[13329] = 12'h1ef;
    rom[13330] = 12'h1ef;
    rom[13331] = 12'h1ef;
    rom[13332] = 12'h1ef;
    rom[13333] = 12'h1ef;
    rom[13334] = 12'h1ef;
    rom[13335] = 12'h1ef;
    rom[13336] = 12'h1ef;
    rom[13337] = 12'h1ef;
    rom[13338] = 12'h1ef;
    rom[13339] = 12'h1ef;
    rom[13340] = 12'h1ef;
    rom[13341] = 12'h1ef;
    rom[13342] = 12'h1ef;
    rom[13343] = 12'h1ee;
    rom[13344] = 12'h1ee;
    rom[13345] = 12'h1ee;
    rom[13346] = 12'h1ee;
    rom[13347] = 12'h1ee;
    rom[13348] = 12'h000;
    rom[13349] = 12'h000;
    rom[13350] = 12'h000;
    rom[13351] = 12'h000;
    rom[13352] = 12'h000;
    rom[13353] = 12'h000;
    rom[13354] = 12'h000;
    rom[13355] = 12'h000;
    rom[13356] = 12'h000;
    rom[13357] = 12'h000;
    rom[13358] = 12'h000;
    rom[13359] = 12'h000;
    rom[13360] = 12'h000;
    rom[13361] = 12'h000;
    rom[13362] = 12'h000;
    rom[13363] = 12'h000;
    rom[13364] = 12'h000;
    rom[13365] = 12'h000;
    rom[13366] = 12'h000;
    rom[13367] = 12'h000;
    rom[13368] = 12'h000;
    rom[13369] = 12'h000;
    rom[13370] = 12'h000;
    rom[13371] = 12'h000;
    rom[13372] = 12'h000;
    rom[13373] = 12'h000;
    rom[13374] = 12'h000;
    rom[13375] = 12'h000;
    rom[13376] = 12'h000;
    rom[13377] = 12'h000;
    rom[13378] = 12'h000;
    rom[13379] = 12'h000;
    rom[13380] = 12'h000;
    rom[13381] = 12'h000;
    rom[13382] = 12'h000;
    rom[13383] = 12'h000;
    rom[13384] = 12'h000;
    rom[13385] = 12'h000;
    rom[13386] = 12'h000;
    rom[13387] = 12'h000;
    rom[13388] = 12'h000;
    rom[13389] = 12'h000;
    rom[13390] = 12'h000;
    rom[13391] = 12'h000;
    rom[13392] = 12'h000;
    rom[13393] = 12'h000;
    rom[13394] = 12'h000;
    rom[13395] = 12'h000;
    rom[13396] = 12'h000;
    rom[13397] = 12'h000;
    rom[13398] = 12'h000;
    rom[13399] = 12'h000;
    rom[13400] = 12'h000;
    rom[13401] = 12'h000;
    rom[13402] = 12'h000;
    rom[13403] = 12'h000;
    rom[13404] = 12'h3a3;
    rom[13405] = 12'h3a3;
    rom[13406] = 12'h3a3;
    rom[13407] = 12'h3a2;
    rom[13408] = 12'h3a2;
    rom[13409] = 12'h3a2;
    rom[13410] = 12'h3a2;
    rom[13411] = 12'h3a2;
    rom[13412] = 12'h3a2;
    rom[13413] = 12'h3a2;
    rom[13414] = 12'h3a2;
    rom[13415] = 12'h3a2;
    rom[13416] = 12'h3a2;
    rom[13417] = 12'h3a2;
    rom[13418] = 12'h3a2;
    rom[13419] = 12'h3a2;
    rom[13420] = 12'h3a2;
    rom[13421] = 12'h3a2;
    rom[13422] = 12'h3a2;
    rom[13423] = 12'h3a2;
    rom[13424] = 12'h3a2;
    rom[13425] = 12'h392;
    rom[13426] = 12'h000;
    rom[13427] = 12'h000;
    rom[13428] = 12'h000;
    rom[13429] = 12'h000;
    rom[13430] = 12'h000;
    rom[13431] = 12'h000;
    rom[13432] = 12'h000;
    rom[13433] = 12'h000;
    rom[13434] = 12'h000;
    rom[13435] = 12'h000;
    rom[13436] = 12'h000;
    rom[13437] = 12'h000;
    rom[13438] = 12'h000;
    rom[13439] = 12'h000;
    rom[13440] = 12'h000;
    rom[13441] = 12'h000;
    rom[13442] = 12'h000;
    rom[13443] = 12'h000;
    rom[13444] = 12'h000;
    rom[13445] = 12'h000;
    rom[13446] = 12'h000;
    rom[13447] = 12'h000;
    rom[13448] = 12'h000;
    rom[13449] = 12'h000;
    rom[13450] = 12'h000;
    rom[13451] = 12'h000;
    rom[13452] = 12'h000;
    rom[13453] = 12'h000;
    rom[13454] = 12'h000;
    rom[13455] = 12'h1ef;
    rom[13456] = 12'h1ef;
    rom[13457] = 12'h1ef;
    rom[13458] = 12'h1ef;
    rom[13459] = 12'h1ef;
    rom[13460] = 12'h1ef;
    rom[13461] = 12'h1ef;
    rom[13462] = 12'h1ef;
    rom[13463] = 12'h1ef;
    rom[13464] = 12'h1ef;
    rom[13465] = 12'h1ef;
    rom[13466] = 12'h1ef;
    rom[13467] = 12'h1ef;
    rom[13468] = 12'h1ef;
    rom[13469] = 12'h1ef;
    rom[13470] = 12'h1ef;
    rom[13471] = 12'h1ee;
    rom[13472] = 12'h1ee;
    rom[13473] = 12'h1ee;
    rom[13474] = 12'h1ee;
    rom[13475] = 12'h1ee;
    rom[13476] = 12'h1ee;
    rom[13477] = 12'h1ee;
    rom[13478] = 12'h000;
    rom[13479] = 12'h000;
    rom[13480] = 12'h000;
    rom[13481] = 12'h000;
    rom[13482] = 12'h000;
    rom[13483] = 12'h000;
    rom[13484] = 12'h000;
    rom[13485] = 12'h000;
    rom[13486] = 12'h000;
    rom[13487] = 12'h000;
    rom[13488] = 12'h000;
    rom[13489] = 12'h000;
    rom[13490] = 12'h000;
    rom[13491] = 12'h000;
    rom[13492] = 12'h000;
    rom[13493] = 12'h000;
    rom[13494] = 12'h000;
    rom[13495] = 12'h000;
    rom[13496] = 12'h000;
    rom[13497] = 12'h000;
    rom[13498] = 12'h000;
    rom[13499] = 12'h000;
    rom[13500] = 12'h000;
    rom[13501] = 12'h000;
    rom[13502] = 12'h000;
    rom[13503] = 12'h000;
    rom[13504] = 12'h000;
    rom[13505] = 12'h000;
    rom[13506] = 12'h000;
    rom[13507] = 12'h000;
    rom[13508] = 12'h000;
    rom[13509] = 12'h000;
    rom[13510] = 12'h000;
    rom[13511] = 12'h000;
    rom[13512] = 12'h000;
    rom[13513] = 12'h000;
    rom[13514] = 12'h000;
    rom[13515] = 12'h000;
    rom[13516] = 12'h000;
    rom[13517] = 12'h000;
    rom[13518] = 12'h000;
    rom[13519] = 12'h000;
    rom[13520] = 12'h000;
    rom[13521] = 12'h000;
    rom[13522] = 12'h000;
    rom[13523] = 12'h000;
    rom[13524] = 12'h000;
    rom[13525] = 12'h000;
    rom[13526] = 12'h000;
    rom[13527] = 12'h000;
    rom[13528] = 12'h000;
    rom[13529] = 12'h000;
    rom[13530] = 12'h3a4;
    rom[13531] = 12'h3a3;
    rom[13532] = 12'h3a3;
    rom[13533] = 12'h3a3;
    rom[13534] = 12'h3a3;
    rom[13535] = 12'h3a2;
    rom[13536] = 12'h3a2;
    rom[13537] = 12'h3a2;
    rom[13538] = 12'h3a2;
    rom[13539] = 12'h3a2;
    rom[13540] = 12'h3a2;
    rom[13541] = 12'h3a2;
    rom[13542] = 12'h3a2;
    rom[13543] = 12'h3a2;
    rom[13544] = 12'h3a2;
    rom[13545] = 12'h3a2;
    rom[13546] = 12'h3a2;
    rom[13547] = 12'h3a2;
    rom[13548] = 12'h3a2;
    rom[13549] = 12'h3a2;
    rom[13550] = 12'h3a2;
    rom[13551] = 12'h3a2;
    rom[13552] = 12'h3a2;
    rom[13553] = 12'h000;
    rom[13554] = 12'h000;
    rom[13555] = 12'h000;
    rom[13556] = 12'h000;
    rom[13557] = 12'h000;
    rom[13558] = 12'h000;
    rom[13559] = 12'h000;
    rom[13560] = 12'h000;
    rom[13561] = 12'h000;
    rom[13562] = 12'h000;
    rom[13563] = 12'h000;
    rom[13564] = 12'h000;
    rom[13565] = 12'h000;
    rom[13566] = 12'h000;
    rom[13567] = 12'h000;
    rom[13568] = 12'h000;
    rom[13569] = 12'h000;
    rom[13570] = 12'h000;
    rom[13571] = 12'h000;
    rom[13572] = 12'h000;
    rom[13573] = 12'h000;
    rom[13574] = 12'h000;
    rom[13575] = 12'h000;
    rom[13576] = 12'h000;
    rom[13577] = 12'h000;
    rom[13578] = 12'h000;
    rom[13579] = 12'h000;
    rom[13580] = 12'h000;
    rom[13581] = 12'h000;
    rom[13582] = 12'h000;
    rom[13583] = 12'h000;
    rom[13584] = 12'h1ef;
    rom[13585] = 12'h1ef;
    rom[13586] = 12'h1ef;
    rom[13587] = 12'h1ef;
    rom[13588] = 12'h1ef;
    rom[13589] = 12'h1ef;
    rom[13590] = 12'h1ef;
    rom[13591] = 12'h1ef;
    rom[13592] = 12'h1ef;
    rom[13593] = 12'h1ef;
    rom[13594] = 12'h1ef;
    rom[13595] = 12'h1ef;
    rom[13596] = 12'h1ef;
    rom[13597] = 12'h1ef;
    rom[13598] = 12'h1ee;
    rom[13599] = 12'h1ee;
    rom[13600] = 12'h1ee;
    rom[13601] = 12'h1ee;
    rom[13602] = 12'h1ee;
    rom[13603] = 12'h1ee;
    rom[13604] = 12'h1ee;
    rom[13605] = 12'h1ee;
    rom[13606] = 12'h1ee;
    rom[13607] = 12'h000;
    rom[13608] = 12'h000;
    rom[13609] = 12'h000;
    rom[13610] = 12'h000;
    rom[13611] = 12'h000;
    rom[13612] = 12'h000;
    rom[13613] = 12'h000;
    rom[13614] = 12'h000;
    rom[13615] = 12'h000;
    rom[13616] = 12'h000;
    rom[13617] = 12'h000;
    rom[13618] = 12'h000;
    rom[13619] = 12'h000;
    rom[13620] = 12'h000;
    rom[13621] = 12'h000;
    rom[13622] = 12'h000;
    rom[13623] = 12'h000;
    rom[13624] = 12'h000;
    rom[13625] = 12'h000;
    rom[13626] = 12'h000;
    rom[13627] = 12'h000;
    rom[13628] = 12'h000;
    rom[13629] = 12'h000;
    rom[13630] = 12'h000;
    rom[13631] = 12'h000;
    rom[13632] = 12'h000;
    rom[13633] = 12'h000;
    rom[13634] = 12'h000;
    rom[13635] = 12'h000;
    rom[13636] = 12'h000;
    rom[13637] = 12'h000;
    rom[13638] = 12'h000;
    rom[13639] = 12'h000;
    rom[13640] = 12'h000;
    rom[13641] = 12'h000;
    rom[13642] = 12'h000;
    rom[13643] = 12'h000;
    rom[13644] = 12'h000;
    rom[13645] = 12'h000;
    rom[13646] = 12'h000;
    rom[13647] = 12'h000;
    rom[13648] = 12'h000;
    rom[13649] = 12'h000;
    rom[13650] = 12'h000;
    rom[13651] = 12'h000;
    rom[13652] = 12'h000;
    rom[13653] = 12'h000;
    rom[13654] = 12'h000;
    rom[13655] = 12'h000;
    rom[13656] = 12'h3b4;
    rom[13657] = 12'h3a4;
    rom[13658] = 12'h3a4;
    rom[13659] = 12'h3a3;
    rom[13660] = 12'h3a3;
    rom[13661] = 12'h3a3;
    rom[13662] = 12'h3a3;
    rom[13663] = 12'h3a2;
    rom[13664] = 12'h3a2;
    rom[13665] = 12'h3a2;
    rom[13666] = 12'h3a2;
    rom[13667] = 12'h3a2;
    rom[13668] = 12'h3a2;
    rom[13669] = 12'h3a2;
    rom[13670] = 12'h3a2;
    rom[13671] = 12'h3a2;
    rom[13672] = 12'h3a2;
    rom[13673] = 12'h3a2;
    rom[13674] = 12'h3a2;
    rom[13675] = 12'h3a2;
    rom[13676] = 12'h3a2;
    rom[13677] = 12'h3a2;
    rom[13678] = 12'h3a2;
    rom[13679] = 12'h3a2;
    rom[13680] = 12'h000;
    rom[13681] = 12'h000;
    rom[13682] = 12'h000;
    rom[13683] = 12'h000;
    rom[13684] = 12'h000;
    rom[13685] = 12'h000;
    rom[13686] = 12'h000;
    rom[13687] = 12'h000;
    rom[13688] = 12'h000;
    rom[13689] = 12'h000;
    rom[13690] = 12'h000;
    rom[13691] = 12'h000;
    rom[13692] = 12'h000;
    rom[13693] = 12'h000;
    rom[13694] = 12'h000;
    rom[13695] = 12'h000;
    rom[13696] = 12'h000;
    rom[13697] = 12'h000;
    rom[13698] = 12'h000;
    rom[13699] = 12'h000;
    rom[13700] = 12'h000;
    rom[13701] = 12'h000;
    rom[13702] = 12'h000;
    rom[13703] = 12'h000;
    rom[13704] = 12'h000;
    rom[13705] = 12'h000;
    rom[13706] = 12'h000;
    rom[13707] = 12'h000;
    rom[13708] = 12'h000;
    rom[13709] = 12'h000;
    rom[13710] = 12'h000;
    rom[13711] = 12'h000;
    rom[13712] = 12'h000;
    rom[13713] = 12'h1ef;
    rom[13714] = 12'h1ef;
    rom[13715] = 12'h1ef;
    rom[13716] = 12'h1ef;
    rom[13717] = 12'h1ef;
    rom[13718] = 12'h1ef;
    rom[13719] = 12'h1ef;
    rom[13720] = 12'h1ef;
    rom[13721] = 12'h1ef;
    rom[13722] = 12'h1ef;
    rom[13723] = 12'h1ef;
    rom[13724] = 12'h1ef;
    rom[13725] = 12'h1ef;
    rom[13726] = 12'h1ee;
    rom[13727] = 12'h1ee;
    rom[13728] = 12'h1ee;
    rom[13729] = 12'h1ee;
    rom[13730] = 12'h1ee;
    rom[13731] = 12'h1ee;
    rom[13732] = 12'h1ee;
    rom[13733] = 12'h1ee;
    rom[13734] = 12'h1ee;
    rom[13735] = 12'h1ee;
    rom[13736] = 12'h1ee;
    rom[13737] = 12'h000;
    rom[13738] = 12'h000;
    rom[13739] = 12'h000;
    rom[13740] = 12'h000;
    rom[13741] = 12'h000;
    rom[13742] = 12'h000;
    rom[13743] = 12'h000;
    rom[13744] = 12'h000;
    rom[13745] = 12'h000;
    rom[13746] = 12'h000;
    rom[13747] = 12'h000;
    rom[13748] = 12'h000;
    rom[13749] = 12'h000;
    rom[13750] = 12'h000;
    rom[13751] = 12'h000;
    rom[13752] = 12'h000;
    rom[13753] = 12'h000;
    rom[13754] = 12'h000;
    rom[13755] = 12'h000;
    rom[13756] = 12'h000;
    rom[13757] = 12'h000;
    rom[13758] = 12'h000;
    rom[13759] = 12'h000;
    rom[13760] = 12'h000;
    rom[13761] = 12'h000;
    rom[13762] = 12'h000;
    rom[13763] = 12'h000;
    rom[13764] = 12'h000;
    rom[13765] = 12'h000;
    rom[13766] = 12'h000;
    rom[13767] = 12'h000;
    rom[13768] = 12'h000;
    rom[13769] = 12'h000;
    rom[13770] = 12'h000;
    rom[13771] = 12'h000;
    rom[13772] = 12'h000;
    rom[13773] = 12'h000;
    rom[13774] = 12'h000;
    rom[13775] = 12'h000;
    rom[13776] = 12'h000;
    rom[13777] = 12'h000;
    rom[13778] = 12'h000;
    rom[13779] = 12'h000;
    rom[13780] = 12'h000;
    rom[13781] = 12'h000;
    rom[13782] = 12'h000;
    rom[13783] = 12'h3a4;
    rom[13784] = 12'h3a4;
    rom[13785] = 12'h3a4;
    rom[13786] = 12'h3a4;
    rom[13787] = 12'h3a3;
    rom[13788] = 12'h3a3;
    rom[13789] = 12'h3a3;
    rom[13790] = 12'h3a3;
    rom[13791] = 12'h3a3;
    rom[13792] = 12'h3a2;
    rom[13793] = 12'h3a2;
    rom[13794] = 12'h3a2;
    rom[13795] = 12'h3a2;
    rom[13796] = 12'h3a2;
    rom[13797] = 12'h3a2;
    rom[13798] = 12'h3a2;
    rom[13799] = 12'h3a2;
    rom[13800] = 12'h3a2;
    rom[13801] = 12'h3a2;
    rom[13802] = 12'h3a2;
    rom[13803] = 12'h3a2;
    rom[13804] = 12'h3a2;
    rom[13805] = 12'h3a2;
    rom[13806] = 12'h3a2;
    rom[13807] = 12'h000;
    rom[13808] = 12'h000;
    rom[13809] = 12'h000;
    rom[13810] = 12'h000;
    rom[13811] = 12'h000;
    rom[13812] = 12'h000;
    rom[13813] = 12'h000;
    rom[13814] = 12'h000;
    rom[13815] = 12'h000;
    rom[13816] = 12'h000;
    rom[13817] = 12'h000;
    rom[13818] = 12'h000;
    rom[13819] = 12'h000;
    rom[13820] = 12'h000;
    rom[13821] = 12'h000;
    rom[13822] = 12'h000;
    rom[13823] = 12'h000;
    rom[13824] = 12'h000;
    rom[13825] = 12'h000;
    rom[13826] = 12'h000;
    rom[13827] = 12'h000;
    rom[13828] = 12'h000;
    rom[13829] = 12'h000;
    rom[13830] = 12'h000;
    rom[13831] = 12'h000;
    rom[13832] = 12'h000;
    rom[13833] = 12'h000;
    rom[13834] = 12'h000;
    rom[13835] = 12'h000;
    rom[13836] = 12'h000;
    rom[13837] = 12'h000;
    rom[13838] = 12'h000;
    rom[13839] = 12'h000;
    rom[13840] = 12'h000;
    rom[13841] = 12'h000;
    rom[13842] = 12'h1ef;
    rom[13843] = 12'h1ef;
    rom[13844] = 12'h1ef;
    rom[13845] = 12'h1ef;
    rom[13846] = 12'h1ef;
    rom[13847] = 12'h1ef;
    rom[13848] = 12'h1ef;
    rom[13849] = 12'h1ef;
    rom[13850] = 12'h1ef;
    rom[13851] = 12'h1ef;
    rom[13852] = 12'h1ef;
    rom[13853] = 12'h1ee;
    rom[13854] = 12'h1ee;
    rom[13855] = 12'h1ee;
    rom[13856] = 12'h1ee;
    rom[13857] = 12'h1ee;
    rom[13858] = 12'h1ee;
    rom[13859] = 12'h1ee;
    rom[13860] = 12'h1ee;
    rom[13861] = 12'h1ee;
    rom[13862] = 12'h1ee;
    rom[13863] = 12'h1ee;
    rom[13864] = 12'h1ee;
    rom[13865] = 12'h1ed;
    rom[13866] = 12'h1ed;
    rom[13867] = 12'h000;
    rom[13868] = 12'h000;
    rom[13869] = 12'h000;
    rom[13870] = 12'h000;
    rom[13871] = 12'h000;
    rom[13872] = 12'h000;
    rom[13873] = 12'h000;
    rom[13874] = 12'h000;
    rom[13875] = 12'h000;
    rom[13876] = 12'h000;
    rom[13877] = 12'h000;
    rom[13878] = 12'h000;
    rom[13879] = 12'h000;
    rom[13880] = 12'h000;
    rom[13881] = 12'h000;
    rom[13882] = 12'h000;
    rom[13883] = 12'h000;
    rom[13884] = 12'h000;
    rom[13885] = 12'h000;
    rom[13886] = 12'h000;
    rom[13887] = 12'h000;
    rom[13888] = 12'h000;
    rom[13889] = 12'h000;
    rom[13890] = 12'h000;
    rom[13891] = 12'h000;
    rom[13892] = 12'h000;
    rom[13893] = 12'h000;
    rom[13894] = 12'h000;
    rom[13895] = 12'h000;
    rom[13896] = 12'h000;
    rom[13897] = 12'h000;
    rom[13898] = 12'h000;
    rom[13899] = 12'h000;
    rom[13900] = 12'h000;
    rom[13901] = 12'h000;
    rom[13902] = 12'h000;
    rom[13903] = 12'h000;
    rom[13904] = 12'h000;
    rom[13905] = 12'h000;
    rom[13906] = 12'h000;
    rom[13907] = 12'h000;
    rom[13908] = 12'h000;
    rom[13909] = 12'h3b5;
    rom[13910] = 12'h3b5;
    rom[13911] = 12'h3a4;
    rom[13912] = 12'h3a4;
    rom[13913] = 12'h3a4;
    rom[13914] = 12'h3a4;
    rom[13915] = 12'h3a3;
    rom[13916] = 12'h3a3;
    rom[13917] = 12'h3a3;
    rom[13918] = 12'h3a3;
    rom[13919] = 12'h3a3;
    rom[13920] = 12'h3a2;
    rom[13921] = 12'h3a2;
    rom[13922] = 12'h3a2;
    rom[13923] = 12'h3a2;
    rom[13924] = 12'h3a2;
    rom[13925] = 12'h3a2;
    rom[13926] = 12'h3a2;
    rom[13927] = 12'h3a2;
    rom[13928] = 12'h3a2;
    rom[13929] = 12'h3a2;
    rom[13930] = 12'h3a2;
    rom[13931] = 12'h3a2;
    rom[13932] = 12'h3a2;
    rom[13933] = 12'h3a2;
    rom[13934] = 12'h000;
    rom[13935] = 12'h000;
    rom[13936] = 12'h000;
    rom[13937] = 12'h000;
    rom[13938] = 12'h000;
    rom[13939] = 12'h000;
    rom[13940] = 12'h000;
    rom[13941] = 12'h000;
    rom[13942] = 12'h000;
    rom[13943] = 12'h000;
    rom[13944] = 12'h000;
    rom[13945] = 12'h000;
    rom[13946] = 12'h000;
    rom[13947] = 12'h000;
    rom[13948] = 12'h000;
    rom[13949] = 12'h000;
    rom[13950] = 12'h000;
    rom[13951] = 12'h000;
    rom[13952] = 12'h000;
    rom[13953] = 12'h000;
    rom[13954] = 12'h000;
    rom[13955] = 12'h000;
    rom[13956] = 12'h000;
    rom[13957] = 12'h000;
    rom[13958] = 12'h000;
    rom[13959] = 12'h000;
    rom[13960] = 12'h000;
    rom[13961] = 12'h000;
    rom[13962] = 12'h000;
    rom[13963] = 12'h000;
    rom[13964] = 12'h000;
    rom[13965] = 12'h000;
    rom[13966] = 12'h000;
    rom[13967] = 12'h000;
    rom[13968] = 12'h000;
    rom[13969] = 12'h000;
    rom[13970] = 12'h000;
    rom[13971] = 12'h1ef;
    rom[13972] = 12'h1ef;
    rom[13973] = 12'h1ef;
    rom[13974] = 12'h1ef;
    rom[13975] = 12'h1ef;
    rom[13976] = 12'h1ef;
    rom[13977] = 12'h1ef;
    rom[13978] = 12'h1ef;
    rom[13979] = 12'h1ef;
    rom[13980] = 12'h1ef;
    rom[13981] = 12'h1ee;
    rom[13982] = 12'h1ee;
    rom[13983] = 12'h1ee;
    rom[13984] = 12'h1ee;
    rom[13985] = 12'h1ee;
    rom[13986] = 12'h1ee;
    rom[13987] = 12'h1ee;
    rom[13988] = 12'h1ee;
    rom[13989] = 12'h1ee;
    rom[13990] = 12'h1ee;
    rom[13991] = 12'h1ee;
    rom[13992] = 12'h1ee;
    rom[13993] = 12'h1ed;
    rom[13994] = 12'h1ed;
    rom[13995] = 12'h1ed;
    rom[13996] = 12'h1ed;
    rom[13997] = 12'h2dd;
    rom[13998] = 12'h000;
    rom[13999] = 12'h000;
    rom[14000] = 12'h000;
    rom[14001] = 12'h000;
    rom[14002] = 12'h000;
    rom[14003] = 12'h000;
    rom[14004] = 12'h000;
    rom[14005] = 12'h000;
    rom[14006] = 12'h000;
    rom[14007] = 12'h000;
    rom[14008] = 12'h000;
    rom[14009] = 12'h000;
    rom[14010] = 12'h000;
    rom[14011] = 12'h000;
    rom[14012] = 12'h000;
    rom[14013] = 12'h000;
    rom[14014] = 12'h000;
    rom[14015] = 12'h000;
    rom[14016] = 12'h000;
    rom[14017] = 12'h000;
    rom[14018] = 12'h000;
    rom[14019] = 12'h000;
    rom[14020] = 12'h000;
    rom[14021] = 12'h000;
    rom[14022] = 12'h000;
    rom[14023] = 12'h000;
    rom[14024] = 12'h000;
    rom[14025] = 12'h000;
    rom[14026] = 12'h000;
    rom[14027] = 12'h000;
    rom[14028] = 12'h000;
    rom[14029] = 12'h000;
    rom[14030] = 12'h000;
    rom[14031] = 12'h000;
    rom[14032] = 12'h000;
    rom[14033] = 12'h000;
    rom[14034] = 12'h3b6;
    rom[14035] = 12'h3b5;
    rom[14036] = 12'h3b5;
    rom[14037] = 12'h3b5;
    rom[14038] = 12'h3b5;
    rom[14039] = 12'h3b4;
    rom[14040] = 12'h3a4;
    rom[14041] = 12'h3a4;
    rom[14042] = 12'h3a4;
    rom[14043] = 12'h3a4;
    rom[14044] = 12'h3a3;
    rom[14045] = 12'h3a3;
    rom[14046] = 12'h3a3;
    rom[14047] = 12'h3a3;
    rom[14048] = 12'h3a2;
    rom[14049] = 12'h3a2;
    rom[14050] = 12'h3a2;
    rom[14051] = 12'h3a2;
    rom[14052] = 12'h3a2;
    rom[14053] = 12'h3a2;
    rom[14054] = 12'h3a2;
    rom[14055] = 12'h3a2;
    rom[14056] = 12'h3a2;
    rom[14057] = 12'h3a2;
    rom[14058] = 12'h3a2;
    rom[14059] = 12'h3a2;
    rom[14060] = 12'h3a2;
    rom[14061] = 12'h000;
    rom[14062] = 12'h000;
    rom[14063] = 12'h000;
    rom[14064] = 12'h000;
    rom[14065] = 12'h000;
    rom[14066] = 12'h000;
    rom[14067] = 12'h000;
    rom[14068] = 12'h000;
    rom[14069] = 12'h000;
    rom[14070] = 12'h000;
    rom[14071] = 12'h000;
    rom[14072] = 12'h000;
    rom[14073] = 12'h000;
    rom[14074] = 12'h000;
    rom[14075] = 12'h000;
    rom[14076] = 12'h000;
    rom[14077] = 12'h000;
    rom[14078] = 12'h000;
    rom[14079] = 12'h000;
    rom[14080] = 12'h000;
    rom[14081] = 12'h000;
    rom[14082] = 12'h000;
    rom[14083] = 12'h000;
    rom[14084] = 12'h000;
    rom[14085] = 12'h000;
    rom[14086] = 12'h000;
    rom[14087] = 12'h000;
    rom[14088] = 12'h000;
    rom[14089] = 12'h000;
    rom[14090] = 12'h000;
    rom[14091] = 12'h000;
    rom[14092] = 12'h000;
    rom[14093] = 12'h000;
    rom[14094] = 12'h000;
    rom[14095] = 12'h000;
    rom[14096] = 12'h000;
    rom[14097] = 12'h000;
    rom[14098] = 12'h000;
    rom[14099] = 12'h000;
    rom[14100] = 12'h1ef;
    rom[14101] = 12'h1ef;
    rom[14102] = 12'h1ef;
    rom[14103] = 12'h1ef;
    rom[14104] = 12'h1ef;
    rom[14105] = 12'h1ef;
    rom[14106] = 12'h1ef;
    rom[14107] = 12'h1ef;
    rom[14108] = 12'h1ef;
    rom[14109] = 12'h1ee;
    rom[14110] = 12'h1ee;
    rom[14111] = 12'h1ee;
    rom[14112] = 12'h1ee;
    rom[14113] = 12'h1ee;
    rom[14114] = 12'h1ee;
    rom[14115] = 12'h1ee;
    rom[14116] = 12'h1ee;
    rom[14117] = 12'h1ee;
    rom[14118] = 12'h1ee;
    rom[14119] = 12'h1ee;
    rom[14120] = 12'h1ed;
    rom[14121] = 12'h1ed;
    rom[14122] = 12'h1ed;
    rom[14123] = 12'h1ed;
    rom[14124] = 12'h1ed;
    rom[14125] = 12'h2dd;
    rom[14126] = 12'h2dd;
    rom[14127] = 12'h2dd;
    rom[14128] = 12'h000;
    rom[14129] = 12'h000;
    rom[14130] = 12'h000;
    rom[14131] = 12'h000;
    rom[14132] = 12'h000;
    rom[14133] = 12'h000;
    rom[14134] = 12'h000;
    rom[14135] = 12'h000;
    rom[14136] = 12'h000;
    rom[14137] = 12'h000;
    rom[14138] = 12'h000;
    rom[14139] = 12'h000;
    rom[14140] = 12'h000;
    rom[14141] = 12'h000;
    rom[14142] = 12'h000;
    rom[14143] = 12'h000;
    rom[14144] = 12'h000;
    rom[14145] = 12'h000;
    rom[14146] = 12'h000;
    rom[14147] = 12'h000;
    rom[14148] = 12'h000;
    rom[14149] = 12'h000;
    rom[14150] = 12'h000;
    rom[14151] = 12'h000;
    rom[14152] = 12'h000;
    rom[14153] = 12'h000;
    rom[14154] = 12'h000;
    rom[14155] = 12'h000;
    rom[14156] = 12'h000;
    rom[14157] = 12'h000;
    rom[14158] = 12'h000;
    rom[14159] = 12'h000;
    rom[14160] = 12'h3b6;
    rom[14161] = 12'h3b6;
    rom[14162] = 12'h3b6;
    rom[14163] = 12'h3b5;
    rom[14164] = 12'h3b5;
    rom[14165] = 12'h3b5;
    rom[14166] = 12'h3b5;
    rom[14167] = 12'h3b4;
    rom[14168] = 12'h3a4;
    rom[14169] = 12'h3a4;
    rom[14170] = 12'h3a4;
    rom[14171] = 12'h3a4;
    rom[14172] = 12'h3a3;
    rom[14173] = 12'h3a3;
    rom[14174] = 12'h3a3;
    rom[14175] = 12'h3a3;
    rom[14176] = 12'h3a2;
    rom[14177] = 12'h3a2;
    rom[14178] = 12'h3a2;
    rom[14179] = 12'h3a2;
    rom[14180] = 12'h3a2;
    rom[14181] = 12'h3a2;
    rom[14182] = 12'h3a2;
    rom[14183] = 12'h3a2;
    rom[14184] = 12'h3a2;
    rom[14185] = 12'h3a2;
    rom[14186] = 12'h3a2;
    rom[14187] = 12'h3a2;
    rom[14188] = 12'h000;
    rom[14189] = 12'h000;
    rom[14190] = 12'h000;
    rom[14191] = 12'h000;
    rom[14192] = 12'h000;
    rom[14193] = 12'h000;
    rom[14194] = 12'h000;
    rom[14195] = 12'h000;
    rom[14196] = 12'h000;
    rom[14197] = 12'h000;
    rom[14198] = 12'h000;
    rom[14199] = 12'h000;
    rom[14200] = 12'h000;
    rom[14201] = 12'h000;
    rom[14202] = 12'h000;
    rom[14203] = 12'h000;
    rom[14204] = 12'h000;
    rom[14205] = 12'h000;
    rom[14206] = 12'h000;
    rom[14207] = 12'h000;
    rom[14208] = 12'h000;
    rom[14209] = 12'h000;
    rom[14210] = 12'h000;
    rom[14211] = 12'h000;
    rom[14212] = 12'h000;
    rom[14213] = 12'h000;
    rom[14214] = 12'h000;
    rom[14215] = 12'h000;
    rom[14216] = 12'h000;
    rom[14217] = 12'h000;
    rom[14218] = 12'h000;
    rom[14219] = 12'h000;
    rom[14220] = 12'h000;
    rom[14221] = 12'h000;
    rom[14222] = 12'h000;
    rom[14223] = 12'h000;
    rom[14224] = 12'h000;
    rom[14225] = 12'h000;
    rom[14226] = 12'h000;
    rom[14227] = 12'h000;
    rom[14228] = 12'h000;
    rom[14229] = 12'h1ef;
    rom[14230] = 12'h1ef;
    rom[14231] = 12'h1ef;
    rom[14232] = 12'h1ef;
    rom[14233] = 12'h1ef;
    rom[14234] = 12'h1ef;
    rom[14235] = 12'h1ef;
    rom[14236] = 12'h1ee;
    rom[14237] = 12'h1ee;
    rom[14238] = 12'h1ee;
    rom[14239] = 12'h1ee;
    rom[14240] = 12'h1ee;
    rom[14241] = 12'h1ee;
    rom[14242] = 12'h1ee;
    rom[14243] = 12'h1ee;
    rom[14244] = 12'h1ee;
    rom[14245] = 12'h1ee;
    rom[14246] = 12'h1ee;
    rom[14247] = 12'h1ee;
    rom[14248] = 12'h1ed;
    rom[14249] = 12'h1ed;
    rom[14250] = 12'h1ed;
    rom[14251] = 12'h1ed;
    rom[14252] = 12'h1ed;
    rom[14253] = 12'h2dd;
    rom[14254] = 12'h2dd;
    rom[14255] = 12'h2dd;
    rom[14256] = 12'h2dc;
    rom[14257] = 12'h2dc;
    rom[14258] = 12'h2dc;
    rom[14259] = 12'h2da;
    rom[14260] = 12'h000;
    rom[14261] = 12'h000;
    rom[14262] = 12'h000;
    rom[14263] = 12'h000;
    rom[14264] = 12'h000;
    rom[14265] = 12'h000;
    rom[14266] = 12'h000;
    rom[14267] = 12'h000;
    rom[14268] = 12'h000;
    rom[14269] = 12'h000;
    rom[14270] = 12'h000;
    rom[14271] = 12'h000;
    rom[14272] = 12'h000;
    rom[14273] = 12'h000;
    rom[14274] = 12'h000;
    rom[14275] = 12'h000;
    rom[14276] = 12'h000;
    rom[14277] = 12'h000;
    rom[14278] = 12'h000;
    rom[14279] = 12'h000;
    rom[14280] = 12'h000;
    rom[14281] = 12'h000;
    rom[14282] = 12'h000;
    rom[14283] = 12'h000;
    rom[14284] = 12'h2b7;
    rom[14285] = 12'h3b7;
    rom[14286] = 12'h3b7;
    rom[14287] = 12'h3b6;
    rom[14288] = 12'h3b6;
    rom[14289] = 12'h3b6;
    rom[14290] = 12'h3b6;
    rom[14291] = 12'h3b5;
    rom[14292] = 12'h3b5;
    rom[14293] = 12'h3b5;
    rom[14294] = 12'h3b5;
    rom[14295] = 12'h3b5;
    rom[14296] = 12'h3a4;
    rom[14297] = 12'h3a4;
    rom[14298] = 12'h3a4;
    rom[14299] = 12'h3a4;
    rom[14300] = 12'h3a3;
    rom[14301] = 12'h3a3;
    rom[14302] = 12'h3a3;
    rom[14303] = 12'h3a3;
    rom[14304] = 12'h3a2;
    rom[14305] = 12'h3a2;
    rom[14306] = 12'h3a2;
    rom[14307] = 12'h3a2;
    rom[14308] = 12'h3a2;
    rom[14309] = 12'h3a2;
    rom[14310] = 12'h3a2;
    rom[14311] = 12'h3a2;
    rom[14312] = 12'h3a2;
    rom[14313] = 12'h3a2;
    rom[14314] = 12'h3a2;
    rom[14315] = 12'h000;
    rom[14316] = 12'h000;
    rom[14317] = 12'h000;
    rom[14318] = 12'h000;
    rom[14319] = 12'h000;
    rom[14320] = 12'h000;
    rom[14321] = 12'h000;
    rom[14322] = 12'h000;
    rom[14323] = 12'h000;
    rom[14324] = 12'h000;
    rom[14325] = 12'h000;
    rom[14326] = 12'h000;
    rom[14327] = 12'h000;
    rom[14328] = 12'h000;
    rom[14329] = 12'h000;
    rom[14330] = 12'h000;
    rom[14331] = 12'h000;
    rom[14332] = 12'h000;
    rom[14333] = 12'h000;
    rom[14334] = 12'h000;
    rom[14335] = 12'h000;
    rom[14336] = 12'h000;
    rom[14337] = 12'h000;
    rom[14338] = 12'h000;
    rom[14339] = 12'h000;
    rom[14340] = 12'h000;
    rom[14341] = 12'h000;
    rom[14342] = 12'h000;
    rom[14343] = 12'h000;
    rom[14344] = 12'h000;
    rom[14345] = 12'h000;
    rom[14346] = 12'h000;
    rom[14347] = 12'h000;
    rom[14348] = 12'h000;
    rom[14349] = 12'h000;
    rom[14350] = 12'h000;
    rom[14351] = 12'h000;
    rom[14352] = 12'h000;
    rom[14353] = 12'h000;
    rom[14354] = 12'h000;
    rom[14355] = 12'h000;
    rom[14356] = 12'h000;
    rom[14357] = 12'h000;
    rom[14358] = 12'h1ef;
    rom[14359] = 12'h1ef;
    rom[14360] = 12'h1ef;
    rom[14361] = 12'h1ef;
    rom[14362] = 12'h1ef;
    rom[14363] = 12'h1ef;
    rom[14364] = 12'h1ee;
    rom[14365] = 12'h1ee;
    rom[14366] = 12'h1ee;
    rom[14367] = 12'h1ee;
    rom[14368] = 12'h1ee;
    rom[14369] = 12'h1ee;
    rom[14370] = 12'h1ee;
    rom[14371] = 12'h1ee;
    rom[14372] = 12'h1ee;
    rom[14373] = 12'h1ee;
    rom[14374] = 12'h1ee;
    rom[14375] = 12'h1ee;
    rom[14376] = 12'h1ed;
    rom[14377] = 12'h1ed;
    rom[14378] = 12'h1ed;
    rom[14379] = 12'h1ed;
    rom[14380] = 12'h2dd;
    rom[14381] = 12'h2dd;
    rom[14382] = 12'h2dd;
    rom[14383] = 12'h2dd;
    rom[14384] = 12'h2dc;
    rom[14385] = 12'h2dc;
    rom[14386] = 12'h2dc;
    rom[14387] = 12'h2dc;
    rom[14388] = 12'h2dc;
    rom[14389] = 12'h2dc;
    rom[14390] = 12'h2db;
    rom[14391] = 12'h2db;
    rom[14392] = 12'h5aa;
    rom[14393] = 12'h000;
    rom[14394] = 12'h000;
    rom[14395] = 12'h000;
    rom[14396] = 12'h000;
    rom[14397] = 12'h000;
    rom[14398] = 12'h000;
    rom[14399] = 12'h000;
    rom[14400] = 12'h000;
    rom[14401] = 12'h000;
    rom[14402] = 12'h000;
    rom[14403] = 12'h000;
    rom[14404] = 12'h000;
    rom[14405] = 12'h000;
    rom[14406] = 12'h000;
    rom[14407] = 12'h2d8;
    rom[14408] = 12'h3c8;
    rom[14409] = 12'h3c8;
    rom[14410] = 12'h3c8;
    rom[14411] = 12'h3c7;
    rom[14412] = 12'h3b7;
    rom[14413] = 12'h3b7;
    rom[14414] = 12'h3b7;
    rom[14415] = 12'h3b6;
    rom[14416] = 12'h3b6;
    rom[14417] = 12'h3b6;
    rom[14418] = 12'h3b6;
    rom[14419] = 12'h3b5;
    rom[14420] = 12'h3b5;
    rom[14421] = 12'h3b5;
    rom[14422] = 12'h3b5;
    rom[14423] = 12'h3b5;
    rom[14424] = 12'h3a4;
    rom[14425] = 12'h3a4;
    rom[14426] = 12'h3a4;
    rom[14427] = 12'h3a4;
    rom[14428] = 12'h3a3;
    rom[14429] = 12'h3a3;
    rom[14430] = 12'h3a3;
    rom[14431] = 12'h3a3;
    rom[14432] = 12'h3a3;
    rom[14433] = 12'h3a2;
    rom[14434] = 12'h3a2;
    rom[14435] = 12'h3a2;
    rom[14436] = 12'h3a2;
    rom[14437] = 12'h3a2;
    rom[14438] = 12'h3a2;
    rom[14439] = 12'h3a2;
    rom[14440] = 12'h3a2;
    rom[14441] = 12'h3a1;
    rom[14442] = 12'h000;
    rom[14443] = 12'h000;
    rom[14444] = 12'h000;
    rom[14445] = 12'h000;
    rom[14446] = 12'h000;
    rom[14447] = 12'h000;
    rom[14448] = 12'h000;
    rom[14449] = 12'h000;
    rom[14450] = 12'h000;
    rom[14451] = 12'h000;
    rom[14452] = 12'h000;
    rom[14453] = 12'h000;
    rom[14454] = 12'h000;
    rom[14455] = 12'h000;
    rom[14456] = 12'h000;
    rom[14457] = 12'h000;
    rom[14458] = 12'h000;
    rom[14459] = 12'h000;
    rom[14460] = 12'h000;
    rom[14461] = 12'h000;
    rom[14462] = 12'h000;
    rom[14463] = 12'h000;
    rom[14464] = 12'h000;
    rom[14465] = 12'h000;
    rom[14466] = 12'h000;
    rom[14467] = 12'h000;
    rom[14468] = 12'h000;
    rom[14469] = 12'h000;
    rom[14470] = 12'h000;
    rom[14471] = 12'h000;
    rom[14472] = 12'h000;
    rom[14473] = 12'h000;
    rom[14474] = 12'h000;
    rom[14475] = 12'h000;
    rom[14476] = 12'h000;
    rom[14477] = 12'h000;
    rom[14478] = 12'h000;
    rom[14479] = 12'h000;
    rom[14480] = 12'h000;
    rom[14481] = 12'h000;
    rom[14482] = 12'h000;
    rom[14483] = 12'h000;
    rom[14484] = 12'h000;
    rom[14485] = 12'h000;
    rom[14486] = 12'h000;
    rom[14487] = 12'h1ef;
    rom[14488] = 12'h1ef;
    rom[14489] = 12'h1ef;
    rom[14490] = 12'h1ef;
    rom[14491] = 12'h1ef;
    rom[14492] = 12'h1ee;
    rom[14493] = 12'h1ee;
    rom[14494] = 12'h1ee;
    rom[14495] = 12'h1ee;
    rom[14496] = 12'h1ee;
    rom[14497] = 12'h1ee;
    rom[14498] = 12'h1ee;
    rom[14499] = 12'h1ee;
    rom[14500] = 12'h1ee;
    rom[14501] = 12'h1ee;
    rom[14502] = 12'h1ee;
    rom[14503] = 12'h1ed;
    rom[14504] = 12'h1ed;
    rom[14505] = 12'h1ed;
    rom[14506] = 12'h1ed;
    rom[14507] = 12'h1ed;
    rom[14508] = 12'h2dd;
    rom[14509] = 12'h2dd;
    rom[14510] = 12'h2dd;
    rom[14511] = 12'h2dc;
    rom[14512] = 12'h2dc;
    rom[14513] = 12'h2dc;
    rom[14514] = 12'h2dc;
    rom[14515] = 12'h2dc;
    rom[14516] = 12'h2dc;
    rom[14517] = 12'h2dc;
    rom[14518] = 12'h2db;
    rom[14519] = 12'h2db;
    rom[14520] = 12'h2db;
    rom[14521] = 12'h2db;
    rom[14522] = 12'h3db;
    rom[14523] = 12'h3db;
    rom[14524] = 12'h3da;
    rom[14525] = 12'h3da;
    rom[14526] = 12'h3ca;
    rom[14527] = 12'h3ca;
    rom[14528] = 12'h3ca;
    rom[14529] = 12'h3ca;
    rom[14530] = 12'h3c9;
    rom[14531] = 12'h3c9;
    rom[14532] = 12'h3c9;
    rom[14533] = 12'h3c9;
    rom[14534] = 12'h3c8;
    rom[14535] = 12'h3c8;
    rom[14536] = 12'h3c8;
    rom[14537] = 12'h3c8;
    rom[14538] = 12'h3c8;
    rom[14539] = 12'h3c7;
    rom[14540] = 12'h3b7;
    rom[14541] = 12'h3b7;
    rom[14542] = 12'h3b7;
    rom[14543] = 12'h3b6;
    rom[14544] = 12'h3b6;
    rom[14545] = 12'h3b6;
    rom[14546] = 12'h3b6;
    rom[14547] = 12'h3b6;
    rom[14548] = 12'h3b5;
    rom[14549] = 12'h3b5;
    rom[14550] = 12'h3b5;
    rom[14551] = 12'h3b5;
    rom[14552] = 12'h3b4;
    rom[14553] = 12'h3a4;
    rom[14554] = 12'h3a4;
    rom[14555] = 12'h3a4;
    rom[14556] = 12'h3a4;
    rom[14557] = 12'h3a3;
    rom[14558] = 12'h3a3;
    rom[14559] = 12'h3a3;
    rom[14560] = 12'h3a3;
    rom[14561] = 12'h3a2;
    rom[14562] = 12'h3a2;
    rom[14563] = 12'h3a2;
    rom[14564] = 12'h3a2;
    rom[14565] = 12'h3a2;
    rom[14566] = 12'h3a2;
    rom[14567] = 12'h3a2;
    rom[14568] = 12'h000;
    rom[14569] = 12'h000;
    rom[14570] = 12'h000;
    rom[14571] = 12'h000;
    rom[14572] = 12'h000;
    rom[14573] = 12'h000;
    rom[14574] = 12'h000;
    rom[14575] = 12'h000;
    rom[14576] = 12'h000;
    rom[14577] = 12'h000;
    rom[14578] = 12'h000;
    rom[14579] = 12'h000;
    rom[14580] = 12'h000;
    rom[14581] = 12'h000;
    rom[14582] = 12'h000;
    rom[14583] = 12'h000;
    rom[14584] = 12'h000;
    rom[14585] = 12'h000;
    rom[14586] = 12'h000;
    rom[14587] = 12'h000;
    rom[14588] = 12'h000;
    rom[14589] = 12'h000;
    rom[14590] = 12'h000;
    rom[14591] = 12'h000;
    rom[14592] = 12'h000;
    rom[14593] = 12'h000;
    rom[14594] = 12'h000;
    rom[14595] = 12'h000;
    rom[14596] = 12'h000;
    rom[14597] = 12'h000;
    rom[14598] = 12'h000;
    rom[14599] = 12'h000;
    rom[14600] = 12'h000;
    rom[14601] = 12'h000;
    rom[14602] = 12'h000;
    rom[14603] = 12'h000;
    rom[14604] = 12'h000;
    rom[14605] = 12'h000;
    rom[14606] = 12'h000;
    rom[14607] = 12'h000;
    rom[14608] = 12'h000;
    rom[14609] = 12'h000;
    rom[14610] = 12'h000;
    rom[14611] = 12'h000;
    rom[14612] = 12'h000;
    rom[14613] = 12'h000;
    rom[14614] = 12'h000;
    rom[14615] = 12'h000;
    rom[14616] = 12'h0ff;
    rom[14617] = 12'h1ef;
    rom[14618] = 12'h1ef;
    rom[14619] = 12'h1ee;
    rom[14620] = 12'h1ee;
    rom[14621] = 12'h1ee;
    rom[14622] = 12'h1ee;
    rom[14623] = 12'h1ee;
    rom[14624] = 12'h1ee;
    rom[14625] = 12'h1ee;
    rom[14626] = 12'h1ee;
    rom[14627] = 12'h1ee;
    rom[14628] = 12'h1ee;
    rom[14629] = 12'h1ee;
    rom[14630] = 12'h1ee;
    rom[14631] = 12'h1ed;
    rom[14632] = 12'h1ed;
    rom[14633] = 12'h1ed;
    rom[14634] = 12'h1ed;
    rom[14635] = 12'h2ed;
    rom[14636] = 12'h2dd;
    rom[14637] = 12'h2dd;
    rom[14638] = 12'h2dd;
    rom[14639] = 12'h2dc;
    rom[14640] = 12'h2dc;
    rom[14641] = 12'h2dc;
    rom[14642] = 12'h2dc;
    rom[14643] = 12'h2dc;
    rom[14644] = 12'h2dc;
    rom[14645] = 12'h2dc;
    rom[14646] = 12'h2db;
    rom[14647] = 12'h2db;
    rom[14648] = 12'h2db;
    rom[14649] = 12'h3db;
    rom[14650] = 12'h3db;
    rom[14651] = 12'h3da;
    rom[14652] = 12'h3da;
    rom[14653] = 12'h3da;
    rom[14654] = 12'h3ca;
    rom[14655] = 12'h3ca;
    rom[14656] = 12'h3ca;
    rom[14657] = 12'h3ca;
    rom[14658] = 12'h3c9;
    rom[14659] = 12'h3c9;
    rom[14660] = 12'h3c9;
    rom[14661] = 12'h3c9;
    rom[14662] = 12'h3c9;
    rom[14663] = 12'h3c8;
    rom[14664] = 12'h3c8;
    rom[14665] = 12'h3c8;
    rom[14666] = 12'h3c8;
    rom[14667] = 12'h3c7;
    rom[14668] = 12'h3b7;
    rom[14669] = 12'h3b7;
    rom[14670] = 12'h3b7;
    rom[14671] = 12'h3b6;
    rom[14672] = 12'h3b6;
    rom[14673] = 12'h3b6;
    rom[14674] = 12'h3b6;
    rom[14675] = 12'h3b6;
    rom[14676] = 12'h3b5;
    rom[14677] = 12'h3b5;
    rom[14678] = 12'h3b5;
    rom[14679] = 12'h3b5;
    rom[14680] = 12'h3b4;
    rom[14681] = 12'h3a4;
    rom[14682] = 12'h3a4;
    rom[14683] = 12'h3a4;
    rom[14684] = 12'h3a4;
    rom[14685] = 12'h3a3;
    rom[14686] = 12'h3a3;
    rom[14687] = 12'h3a3;
    rom[14688] = 12'h3a3;
    rom[14689] = 12'h3a2;
    rom[14690] = 12'h3a2;
    rom[14691] = 12'h3a2;
    rom[14692] = 12'h3a2;
    rom[14693] = 12'h3a2;
    rom[14694] = 12'h3a2;
    rom[14695] = 12'h000;
    rom[14696] = 12'h000;
    rom[14697] = 12'h000;
    rom[14698] = 12'h000;
    rom[14699] = 12'h000;
    rom[14700] = 12'h000;
    rom[14701] = 12'h000;
    rom[14702] = 12'h000;
    rom[14703] = 12'h000;
    rom[14704] = 12'h000;
    rom[14705] = 12'h000;
    rom[14706] = 12'h000;
    rom[14707] = 12'h000;
    rom[14708] = 12'h000;
    rom[14709] = 12'h000;
    rom[14710] = 12'h000;
    rom[14711] = 12'h000;
    rom[14712] = 12'h000;
    rom[14713] = 12'h000;
    rom[14714] = 12'h000;
    rom[14715] = 12'h000;
    rom[14716] = 12'h000;
    rom[14717] = 12'h000;
    rom[14718] = 12'h000;
    rom[14719] = 12'h000;
    rom[14720] = 12'h000;
    rom[14721] = 12'h000;
    rom[14722] = 12'h000;
    rom[14723] = 12'h000;
    rom[14724] = 12'h000;
    rom[14725] = 12'h000;
    rom[14726] = 12'h000;
    rom[14727] = 12'h000;
    rom[14728] = 12'h000;
    rom[14729] = 12'h000;
    rom[14730] = 12'h000;
    rom[14731] = 12'h000;
    rom[14732] = 12'h000;
    rom[14733] = 12'h000;
    rom[14734] = 12'h000;
    rom[14735] = 12'h000;
    rom[14736] = 12'h000;
    rom[14737] = 12'h000;
    rom[14738] = 12'h000;
    rom[14739] = 12'h000;
    rom[14740] = 12'h000;
    rom[14741] = 12'h000;
    rom[14742] = 12'h000;
    rom[14743] = 12'h000;
    rom[14744] = 12'h000;
    rom[14745] = 12'h000;
    rom[14746] = 12'h1ef;
    rom[14747] = 12'h1ee;
    rom[14748] = 12'h1ee;
    rom[14749] = 12'h1ee;
    rom[14750] = 12'h1ee;
    rom[14751] = 12'h1ee;
    rom[14752] = 12'h1ee;
    rom[14753] = 12'h1ee;
    rom[14754] = 12'h1ee;
    rom[14755] = 12'h1ee;
    rom[14756] = 12'h1ee;
    rom[14757] = 12'h1ee;
    rom[14758] = 12'h1ee;
    rom[14759] = 12'h1ed;
    rom[14760] = 12'h1ed;
    rom[14761] = 12'h1ed;
    rom[14762] = 12'h1ed;
    rom[14763] = 12'h2dd;
    rom[14764] = 12'h2dd;
    rom[14765] = 12'h2dd;
    rom[14766] = 12'h2dc;
    rom[14767] = 12'h2dc;
    rom[14768] = 12'h2dc;
    rom[14769] = 12'h2dc;
    rom[14770] = 12'h2dc;
    rom[14771] = 12'h2dc;
    rom[14772] = 12'h2dc;
    rom[14773] = 12'h2db;
    rom[14774] = 12'h2db;
    rom[14775] = 12'h2db;
    rom[14776] = 12'h2db;
    rom[14777] = 12'h3db;
    rom[14778] = 12'h3db;
    rom[14779] = 12'h3da;
    rom[14780] = 12'h3da;
    rom[14781] = 12'h3ca;
    rom[14782] = 12'h3ca;
    rom[14783] = 12'h3ca;
    rom[14784] = 12'h3ca;
    rom[14785] = 12'h3ca;
    rom[14786] = 12'h3ca;
    rom[14787] = 12'h3c9;
    rom[14788] = 12'h3c9;
    rom[14789] = 12'h3c9;
    rom[14790] = 12'h3c9;
    rom[14791] = 12'h3c8;
    rom[14792] = 12'h3c8;
    rom[14793] = 12'h3c8;
    rom[14794] = 12'h3c8;
    rom[14795] = 12'h3c7;
    rom[14796] = 12'h3b7;
    rom[14797] = 12'h3b7;
    rom[14798] = 12'h3b7;
    rom[14799] = 12'h3b7;
    rom[14800] = 12'h3b6;
    rom[14801] = 12'h3b6;
    rom[14802] = 12'h3b6;
    rom[14803] = 12'h3b6;
    rom[14804] = 12'h3b5;
    rom[14805] = 12'h3b5;
    rom[14806] = 12'h3b5;
    rom[14807] = 12'h3b5;
    rom[14808] = 12'h3b5;
    rom[14809] = 12'h3a4;
    rom[14810] = 12'h3a4;
    rom[14811] = 12'h3a4;
    rom[14812] = 12'h3a4;
    rom[14813] = 12'h3a3;
    rom[14814] = 12'h3a3;
    rom[14815] = 12'h3a3;
    rom[14816] = 12'h3a3;
    rom[14817] = 12'h3a2;
    rom[14818] = 12'h3a2;
    rom[14819] = 12'h3a2;
    rom[14820] = 12'h3a2;
    rom[14821] = 12'h3a2;
    rom[14822] = 12'h000;
    rom[14823] = 12'h000;
    rom[14824] = 12'h000;
    rom[14825] = 12'h000;
    rom[14826] = 12'h000;
    rom[14827] = 12'h000;
    rom[14828] = 12'h000;
    rom[14829] = 12'h000;
    rom[14830] = 12'h000;
    rom[14831] = 12'h000;
    rom[14832] = 12'h000;
    rom[14833] = 12'h000;
    rom[14834] = 12'h000;
    rom[14835] = 12'h000;
    rom[14836] = 12'h000;
    rom[14837] = 12'h000;
    rom[14838] = 12'h000;
    rom[14839] = 12'h000;
    rom[14840] = 12'h000;
    rom[14841] = 12'h000;
    rom[14842] = 12'h000;
    rom[14843] = 12'h000;
    rom[14844] = 12'h000;
    rom[14845] = 12'h000;
    rom[14846] = 12'h000;
    rom[14847] = 12'h000;
    rom[14848] = 12'h000;
    rom[14849] = 12'h000;
    rom[14850] = 12'h000;
    rom[14851] = 12'h000;
    rom[14852] = 12'h000;
    rom[14853] = 12'h000;
    rom[14854] = 12'h000;
    rom[14855] = 12'h000;
    rom[14856] = 12'h000;
    rom[14857] = 12'h000;
    rom[14858] = 12'h000;
    rom[14859] = 12'h000;
    rom[14860] = 12'h000;
    rom[14861] = 12'h000;
    rom[14862] = 12'h000;
    rom[14863] = 12'h000;
    rom[14864] = 12'h000;
    rom[14865] = 12'h000;
    rom[14866] = 12'h000;
    rom[14867] = 12'h000;
    rom[14868] = 12'h000;
    rom[14869] = 12'h000;
    rom[14870] = 12'h000;
    rom[14871] = 12'h000;
    rom[14872] = 12'h000;
    rom[14873] = 12'h000;
    rom[14874] = 12'h000;
    rom[14875] = 12'h1ee;
    rom[14876] = 12'h1ee;
    rom[14877] = 12'h1ee;
    rom[14878] = 12'h1ee;
    rom[14879] = 12'h1ee;
    rom[14880] = 12'h1ee;
    rom[14881] = 12'h1ee;
    rom[14882] = 12'h1ee;
    rom[14883] = 12'h1ee;
    rom[14884] = 12'h1ee;
    rom[14885] = 12'h1ee;
    rom[14886] = 12'h1ed;
    rom[14887] = 12'h1ed;
    rom[14888] = 12'h1ed;
    rom[14889] = 12'h1ed;
    rom[14890] = 12'h1ed;
    rom[14891] = 12'h2dd;
    rom[14892] = 12'h2dd;
    rom[14893] = 12'h2dd;
    rom[14894] = 12'h2dc;
    rom[14895] = 12'h2dc;
    rom[14896] = 12'h2dc;
    rom[14897] = 12'h2dc;
    rom[14898] = 12'h2dc;
    rom[14899] = 12'h2dc;
    rom[14900] = 12'h2dc;
    rom[14901] = 12'h2db;
    rom[14902] = 12'h2db;
    rom[14903] = 12'h2db;
    rom[14904] = 12'h3db;
    rom[14905] = 12'h3db;
    rom[14906] = 12'h3db;
    rom[14907] = 12'h3da;
    rom[14908] = 12'h3da;
    rom[14909] = 12'h3ca;
    rom[14910] = 12'h3ca;
    rom[14911] = 12'h3ca;
    rom[14912] = 12'h3ca;
    rom[14913] = 12'h3ca;
    rom[14914] = 12'h3ca;
    rom[14915] = 12'h3c9;
    rom[14916] = 12'h3c9;
    rom[14917] = 12'h3c9;
    rom[14918] = 12'h3c9;
    rom[14919] = 12'h3c8;
    rom[14920] = 12'h3c8;
    rom[14921] = 12'h3c8;
    rom[14922] = 12'h3c8;
    rom[14923] = 12'h3c7;
    rom[14924] = 12'h3c7;
    rom[14925] = 12'h3b7;
    rom[14926] = 12'h3b7;
    rom[14927] = 12'h3b7;
    rom[14928] = 12'h3b6;
    rom[14929] = 12'h3b6;
    rom[14930] = 12'h3b6;
    rom[14931] = 12'h3b6;
    rom[14932] = 12'h3b5;
    rom[14933] = 12'h3b5;
    rom[14934] = 12'h3b5;
    rom[14935] = 12'h3b5;
    rom[14936] = 12'h3b5;
    rom[14937] = 12'h3a4;
    rom[14938] = 12'h3a4;
    rom[14939] = 12'h3a4;
    rom[14940] = 12'h3a4;
    rom[14941] = 12'h3a3;
    rom[14942] = 12'h3a3;
    rom[14943] = 12'h3a3;
    rom[14944] = 12'h3a3;
    rom[14945] = 12'h3a3;
    rom[14946] = 12'h3a2;
    rom[14947] = 12'h3a2;
    rom[14948] = 12'h000;
    rom[14949] = 12'h000;
    rom[14950] = 12'h000;
    rom[14951] = 12'h000;
    rom[14952] = 12'h000;
    rom[14953] = 12'h000;
    rom[14954] = 12'h000;
    rom[14955] = 12'h000;
    rom[14956] = 12'h000;
    rom[14957] = 12'h000;
    rom[14958] = 12'h000;
    rom[14959] = 12'h000;
    rom[14960] = 12'h000;
    rom[14961] = 12'h000;
    rom[14962] = 12'h000;
    rom[14963] = 12'h000;
    rom[14964] = 12'h000;
    rom[14965] = 12'h000;
    rom[14966] = 12'h000;
    rom[14967] = 12'h000;
    rom[14968] = 12'h000;
    rom[14969] = 12'h000;
    rom[14970] = 12'h000;
    rom[14971] = 12'h000;
    rom[14972] = 12'h000;
    rom[14973] = 12'h000;
    rom[14974] = 12'h000;
    rom[14975] = 12'h000;
    rom[14976] = 12'h000;
    rom[14977] = 12'h000;
    rom[14978] = 12'h000;
    rom[14979] = 12'h000;
    rom[14980] = 12'h000;
    rom[14981] = 12'h000;
    rom[14982] = 12'h000;
    rom[14983] = 12'h000;
    rom[14984] = 12'h000;
    rom[14985] = 12'h000;
    rom[14986] = 12'h000;
    rom[14987] = 12'h000;
    rom[14988] = 12'h000;
    rom[14989] = 12'h000;
    rom[14990] = 12'h000;
    rom[14991] = 12'h000;
    rom[14992] = 12'h000;
    rom[14993] = 12'h000;
    rom[14994] = 12'h000;
    rom[14995] = 12'h000;
    rom[14996] = 12'h000;
    rom[14997] = 12'h000;
    rom[14998] = 12'h000;
    rom[14999] = 12'h000;
    rom[15000] = 12'h000;
    rom[15001] = 12'h000;
    rom[15002] = 12'h000;
    rom[15003] = 12'h000;
    rom[15004] = 12'h000;
    rom[15005] = 12'h1ee;
    rom[15006] = 12'h1ee;
    rom[15007] = 12'h1ee;
    rom[15008] = 12'h1ee;
    rom[15009] = 12'h1ee;
    rom[15010] = 12'h1ee;
    rom[15011] = 12'h1ee;
    rom[15012] = 12'h1ee;
    rom[15013] = 12'h1ee;
    rom[15014] = 12'h1ed;
    rom[15015] = 12'h1ed;
    rom[15016] = 12'h1ed;
    rom[15017] = 12'h1ed;
    rom[15018] = 12'h2dd;
    rom[15019] = 12'h2dd;
    rom[15020] = 12'h2dd;
    rom[15021] = 12'h2dd;
    rom[15022] = 12'h2dc;
    rom[15023] = 12'h2dc;
    rom[15024] = 12'h2dc;
    rom[15025] = 12'h2dc;
    rom[15026] = 12'h2dc;
    rom[15027] = 12'h2dc;
    rom[15028] = 12'h2db;
    rom[15029] = 12'h2db;
    rom[15030] = 12'h2db;
    rom[15031] = 12'h2db;
    rom[15032] = 12'h3db;
    rom[15033] = 12'h3db;
    rom[15034] = 12'h3da;
    rom[15035] = 12'h3da;
    rom[15036] = 12'h3ca;
    rom[15037] = 12'h3ca;
    rom[15038] = 12'h3ca;
    rom[15039] = 12'h3ca;
    rom[15040] = 12'h3ca;
    rom[15041] = 12'h3ca;
    rom[15042] = 12'h3ca;
    rom[15043] = 12'h3c9;
    rom[15044] = 12'h3c9;
    rom[15045] = 12'h3c9;
    rom[15046] = 12'h3c9;
    rom[15047] = 12'h3c8;
    rom[15048] = 12'h3c8;
    rom[15049] = 12'h3c8;
    rom[15050] = 12'h3c8;
    rom[15051] = 12'h3c8;
    rom[15052] = 12'h3c7;
    rom[15053] = 12'h3b7;
    rom[15054] = 12'h3b7;
    rom[15055] = 12'h3b7;
    rom[15056] = 12'h3b6;
    rom[15057] = 12'h3b6;
    rom[15058] = 12'h3b6;
    rom[15059] = 12'h3b6;
    rom[15060] = 12'h3b6;
    rom[15061] = 12'h3b5;
    rom[15062] = 12'h3b5;
    rom[15063] = 12'h3b5;
    rom[15064] = 12'h3b5;
    rom[15065] = 12'h3b4;
    rom[15066] = 12'h3a4;
    rom[15067] = 12'h3a4;
    rom[15068] = 12'h3a4;
    rom[15069] = 12'h3a3;
    rom[15070] = 12'h3a3;
    rom[15071] = 12'h3a3;
    rom[15072] = 12'h3a3;
    rom[15073] = 12'h3a3;
    rom[15074] = 12'h3a2;
    rom[15075] = 12'h000;
    rom[15076] = 12'h000;
    rom[15077] = 12'h000;
    rom[15078] = 12'h000;
    rom[15079] = 12'h000;
    rom[15080] = 12'h000;
    rom[15081] = 12'h000;
    rom[15082] = 12'h000;
    rom[15083] = 12'h000;
    rom[15084] = 12'h000;
    rom[15085] = 12'h000;
    rom[15086] = 12'h000;
    rom[15087] = 12'h000;
    rom[15088] = 12'h000;
    rom[15089] = 12'h000;
    rom[15090] = 12'h000;
    rom[15091] = 12'h000;
    rom[15092] = 12'h000;
    rom[15093] = 12'h000;
    rom[15094] = 12'h000;
    rom[15095] = 12'h000;
    rom[15096] = 12'h000;
    rom[15097] = 12'h000;
    rom[15098] = 12'h000;
    rom[15099] = 12'h000;
    rom[15100] = 12'h000;
    rom[15101] = 12'h000;
    rom[15102] = 12'h000;
    rom[15103] = 12'h000;
    rom[15104] = 12'h000;
    rom[15105] = 12'h000;
    rom[15106] = 12'h000;
    rom[15107] = 12'h000;
    rom[15108] = 12'h000;
    rom[15109] = 12'h000;
    rom[15110] = 12'h000;
    rom[15111] = 12'h000;
    rom[15112] = 12'h000;
    rom[15113] = 12'h000;
    rom[15114] = 12'h000;
    rom[15115] = 12'h000;
    rom[15116] = 12'h000;
    rom[15117] = 12'h000;
    rom[15118] = 12'h000;
    rom[15119] = 12'h000;
    rom[15120] = 12'h000;
    rom[15121] = 12'h000;
    rom[15122] = 12'h000;
    rom[15123] = 12'h000;
    rom[15124] = 12'h000;
    rom[15125] = 12'h000;
    rom[15126] = 12'h000;
    rom[15127] = 12'h000;
    rom[15128] = 12'h000;
    rom[15129] = 12'h000;
    rom[15130] = 12'h000;
    rom[15131] = 12'h000;
    rom[15132] = 12'h000;
    rom[15133] = 12'h000;
    rom[15134] = 12'h1ee;
    rom[15135] = 12'h1ee;
    rom[15136] = 12'h1ee;
    rom[15137] = 12'h1ee;
    rom[15138] = 12'h1ee;
    rom[15139] = 12'h1ee;
    rom[15140] = 12'h1ee;
    rom[15141] = 12'h1ee;
    rom[15142] = 12'h1ed;
    rom[15143] = 12'h1ed;
    rom[15144] = 12'h1ed;
    rom[15145] = 12'h1ed;
    rom[15146] = 12'h2dd;
    rom[15147] = 12'h2dd;
    rom[15148] = 12'h2dd;
    rom[15149] = 12'h2dc;
    rom[15150] = 12'h2dc;
    rom[15151] = 12'h2dc;
    rom[15152] = 12'h2dc;
    rom[15153] = 12'h2dc;
    rom[15154] = 12'h2dc;
    rom[15155] = 12'h2dc;
    rom[15156] = 12'h2db;
    rom[15157] = 12'h2db;
    rom[15158] = 12'h2db;
    rom[15159] = 12'h2db;
    rom[15160] = 12'h3db;
    rom[15161] = 12'h3db;
    rom[15162] = 12'h3da;
    rom[15163] = 12'h3da;
    rom[15164] = 12'h3ca;
    rom[15165] = 12'h3ca;
    rom[15166] = 12'h3ca;
    rom[15167] = 12'h3ca;
    rom[15168] = 12'h3ca;
    rom[15169] = 12'h3ca;
    rom[15170] = 12'h3ca;
    rom[15171] = 12'h3c9;
    rom[15172] = 12'h3c9;
    rom[15173] = 12'h3c9;
    rom[15174] = 12'h3c9;
    rom[15175] = 12'h3c9;
    rom[15176] = 12'h3c8;
    rom[15177] = 12'h3c8;
    rom[15178] = 12'h3c8;
    rom[15179] = 12'h3c8;
    rom[15180] = 12'h3c7;
    rom[15181] = 12'h3b7;
    rom[15182] = 12'h3b7;
    rom[15183] = 12'h3b7;
    rom[15184] = 12'h3b6;
    rom[15185] = 12'h3b6;
    rom[15186] = 12'h3b6;
    rom[15187] = 12'h3b6;
    rom[15188] = 12'h3b6;
    rom[15189] = 12'h3b5;
    rom[15190] = 12'h3b5;
    rom[15191] = 12'h3b5;
    rom[15192] = 12'h3b5;
    rom[15193] = 12'h3b4;
    rom[15194] = 12'h3a4;
    rom[15195] = 12'h3a4;
    rom[15196] = 12'h3a4;
    rom[15197] = 12'h3a4;
    rom[15198] = 12'h3a3;
    rom[15199] = 12'h3a3;
    rom[15200] = 12'h3a3;
    rom[15201] = 12'h000;
    rom[15202] = 12'h000;
    rom[15203] = 12'h000;
    rom[15204] = 12'h000;
    rom[15205] = 12'h000;
    rom[15206] = 12'h000;
    rom[15207] = 12'h000;
    rom[15208] = 12'h000;
    rom[15209] = 12'h000;
    rom[15210] = 12'h000;
    rom[15211] = 12'h000;
    rom[15212] = 12'h000;
    rom[15213] = 12'h000;
    rom[15214] = 12'h000;
    rom[15215] = 12'h000;
    rom[15216] = 12'h000;
    rom[15217] = 12'h000;
    rom[15218] = 12'h000;
    rom[15219] = 12'h000;
    rom[15220] = 12'h000;
    rom[15221] = 12'h000;
    rom[15222] = 12'h000;
    rom[15223] = 12'h000;
    rom[15224] = 12'h000;
    rom[15225] = 12'h000;
    rom[15226] = 12'h000;
    rom[15227] = 12'h000;
    rom[15228] = 12'h000;
    rom[15229] = 12'h000;
    rom[15230] = 12'h000;
    rom[15231] = 12'h000;
    rom[15232] = 12'h000;
    rom[15233] = 12'h000;
    rom[15234] = 12'h000;
    rom[15235] = 12'h000;
    rom[15236] = 12'h000;
    rom[15237] = 12'h000;
    rom[15238] = 12'h000;
    rom[15239] = 12'h000;
    rom[15240] = 12'h000;
    rom[15241] = 12'h000;
    rom[15242] = 12'h000;
    rom[15243] = 12'h000;
    rom[15244] = 12'h000;
    rom[15245] = 12'h000;
    rom[15246] = 12'h000;
    rom[15247] = 12'h000;
    rom[15248] = 12'h000;
    rom[15249] = 12'h000;
    rom[15250] = 12'h000;
    rom[15251] = 12'h000;
    rom[15252] = 12'h000;
    rom[15253] = 12'h000;
    rom[15254] = 12'h000;
    rom[15255] = 12'h000;
    rom[15256] = 12'h000;
    rom[15257] = 12'h000;
    rom[15258] = 12'h000;
    rom[15259] = 12'h000;
    rom[15260] = 12'h000;
    rom[15261] = 12'h000;
    rom[15262] = 12'h000;
    rom[15263] = 12'h000;
    rom[15264] = 12'h1ee;
    rom[15265] = 12'h1ee;
    rom[15266] = 12'h1ee;
    rom[15267] = 12'h1ee;
    rom[15268] = 12'h1ee;
    rom[15269] = 12'h1ed;
    rom[15270] = 12'h1ed;
    rom[15271] = 12'h1ed;
    rom[15272] = 12'h1ed;
    rom[15273] = 12'h2ed;
    rom[15274] = 12'h2dd;
    rom[15275] = 12'h2dd;
    rom[15276] = 12'h2dd;
    rom[15277] = 12'h2dc;
    rom[15278] = 12'h2dc;
    rom[15279] = 12'h2dc;
    rom[15280] = 12'h2dc;
    rom[15281] = 12'h2dc;
    rom[15282] = 12'h2dc;
    rom[15283] = 12'h2dc;
    rom[15284] = 12'h2db;
    rom[15285] = 12'h2db;
    rom[15286] = 12'h2db;
    rom[15287] = 12'h3db;
    rom[15288] = 12'h3db;
    rom[15289] = 12'h3db;
    rom[15290] = 12'h3da;
    rom[15291] = 12'h3da;
    rom[15292] = 12'h3ca;
    rom[15293] = 12'h3ca;
    rom[15294] = 12'h3ca;
    rom[15295] = 12'h3ca;
    rom[15296] = 12'h3ca;
    rom[15297] = 12'h3ca;
    rom[15298] = 12'h3ca;
    rom[15299] = 12'h3ca;
    rom[15300] = 12'h3c9;
    rom[15301] = 12'h3c9;
    rom[15302] = 12'h3c9;
    rom[15303] = 12'h3c9;
    rom[15304] = 12'h3c8;
    rom[15305] = 12'h3c8;
    rom[15306] = 12'h3c8;
    rom[15307] = 12'h3c8;
    rom[15308] = 12'h3c7;
    rom[15309] = 12'h3b7;
    rom[15310] = 12'h3b7;
    rom[15311] = 12'h3b7;
    rom[15312] = 12'h3b7;
    rom[15313] = 12'h3b6;
    rom[15314] = 12'h3b6;
    rom[15315] = 12'h3b6;
    rom[15316] = 12'h3b6;
    rom[15317] = 12'h3b5;
    rom[15318] = 12'h3b5;
    rom[15319] = 12'h3b5;
    rom[15320] = 12'h3b5;
    rom[15321] = 12'h3b4;
    rom[15322] = 12'h3a4;
    rom[15323] = 12'h3a4;
    rom[15324] = 12'h3a4;
    rom[15325] = 12'h3a4;
    rom[15326] = 12'h3a3;
    rom[15327] = 12'h3a3;
    rom[15328] = 12'h000;
    rom[15329] = 12'h000;
    rom[15330] = 12'h000;
    rom[15331] = 12'h000;
    rom[15332] = 12'h000;
    rom[15333] = 12'h000;
    rom[15334] = 12'h000;
    rom[15335] = 12'h000;
    rom[15336] = 12'h000;
    rom[15337] = 12'h000;
    rom[15338] = 12'h000;
    rom[15339] = 12'h000;
    rom[15340] = 12'h000;
    rom[15341] = 12'h000;
    rom[15342] = 12'h000;
    rom[15343] = 12'h000;
    rom[15344] = 12'h000;
    rom[15345] = 12'h000;
    rom[15346] = 12'h000;
    rom[15347] = 12'h000;
    rom[15348] = 12'h000;
    rom[15349] = 12'h000;
    rom[15350] = 12'h000;
    rom[15351] = 12'h000;
    rom[15352] = 12'h000;
    rom[15353] = 12'h000;
    rom[15354] = 12'h000;
    rom[15355] = 12'h000;
    rom[15356] = 12'h000;
    rom[15357] = 12'h000;
    rom[15358] = 12'h000;
    rom[15359] = 12'h000;
    rom[15360] = 12'h000;
    rom[15361] = 12'h000;
    rom[15362] = 12'h000;
    rom[15363] = 12'h000;
    rom[15364] = 12'h000;
    rom[15365] = 12'h000;
    rom[15366] = 12'h000;
    rom[15367] = 12'h000;
    rom[15368] = 12'h000;
    rom[15369] = 12'h000;
    rom[15370] = 12'h000;
    rom[15371] = 12'h000;
    rom[15372] = 12'h000;
    rom[15373] = 12'h000;
    rom[15374] = 12'h000;
    rom[15375] = 12'h000;
    rom[15376] = 12'h000;
    rom[15377] = 12'h000;
    rom[15378] = 12'h000;
    rom[15379] = 12'h000;
    rom[15380] = 12'h000;
    rom[15381] = 12'h000;
    rom[15382] = 12'h000;
    rom[15383] = 12'h000;
    rom[15384] = 12'h000;
    rom[15385] = 12'h000;
    rom[15386] = 12'h000;
    rom[15387] = 12'h000;
    rom[15388] = 12'h000;
    rom[15389] = 12'h000;
    rom[15390] = 12'h000;
    rom[15391] = 12'h000;
    rom[15392] = 12'h000;
    rom[15393] = 12'h000;
    rom[15394] = 12'h1ee;
    rom[15395] = 12'h1ee;
    rom[15396] = 12'h1ee;
    rom[15397] = 12'h1ed;
    rom[15398] = 12'h1ed;
    rom[15399] = 12'h1ed;
    rom[15400] = 12'h1ed;
    rom[15401] = 12'h2dd;
    rom[15402] = 12'h2dd;
    rom[15403] = 12'h2dd;
    rom[15404] = 12'h2dd;
    rom[15405] = 12'h2dc;
    rom[15406] = 12'h2dc;
    rom[15407] = 12'h2dc;
    rom[15408] = 12'h2dc;
    rom[15409] = 12'h2dc;
    rom[15410] = 12'h2dc;
    rom[15411] = 12'h2db;
    rom[15412] = 12'h2db;
    rom[15413] = 12'h2db;
    rom[15414] = 12'h2db;
    rom[15415] = 12'h3db;
    rom[15416] = 12'h3db;
    rom[15417] = 12'h3da;
    rom[15418] = 12'h3da;
    rom[15419] = 12'h3ca;
    rom[15420] = 12'h3ca;
    rom[15421] = 12'h3ca;
    rom[15422] = 12'h3ca;
    rom[15423] = 12'h3ca;
    rom[15424] = 12'h3ca;
    rom[15425] = 12'h3ca;
    rom[15426] = 12'h3ca;
    rom[15427] = 12'h3ca;
    rom[15428] = 12'h3c9;
    rom[15429] = 12'h3c9;
    rom[15430] = 12'h3c9;
    rom[15431] = 12'h3c9;
    rom[15432] = 12'h3c8;
    rom[15433] = 12'h3c8;
    rom[15434] = 12'h3c8;
    rom[15435] = 12'h3c8;
    rom[15436] = 12'h3c7;
    rom[15437] = 12'h3b7;
    rom[15438] = 12'h3b7;
    rom[15439] = 12'h3b7;
    rom[15440] = 12'h3b7;
    rom[15441] = 12'h3b6;
    rom[15442] = 12'h3b6;
    rom[15443] = 12'h3b6;
    rom[15444] = 12'h3b6;
    rom[15445] = 12'h3b5;
    rom[15446] = 12'h3b5;
    rom[15447] = 12'h3b5;
    rom[15448] = 12'h3b5;
    rom[15449] = 12'h3b5;
    rom[15450] = 12'h3a4;
    rom[15451] = 12'h3a4;
    rom[15452] = 12'h3a4;
    rom[15453] = 12'h3a4;
    rom[15454] = 12'h000;
    rom[15455] = 12'h000;
    rom[15456] = 12'h000;
    rom[15457] = 12'h000;
    rom[15458] = 12'h000;
    rom[15459] = 12'h000;
    rom[15460] = 12'h000;
    rom[15461] = 12'h000;
    rom[15462] = 12'h000;
    rom[15463] = 12'h000;
    rom[15464] = 12'h000;
    rom[15465] = 12'h000;
    rom[15466] = 12'h000;
    rom[15467] = 12'h000;
    rom[15468] = 12'h000;
    rom[15469] = 12'h000;
    rom[15470] = 12'h000;
    rom[15471] = 12'h000;
    rom[15472] = 12'h000;
    rom[15473] = 12'h000;
    rom[15474] = 12'h000;
    rom[15475] = 12'h000;
    rom[15476] = 12'h000;
    rom[15477] = 12'h000;
    rom[15478] = 12'h000;
    rom[15479] = 12'h000;
    rom[15480] = 12'h000;
    rom[15481] = 12'h000;
    rom[15482] = 12'h000;
    rom[15483] = 12'h000;
    rom[15484] = 12'h000;
    rom[15485] = 12'h000;
    rom[15486] = 12'h000;
    rom[15487] = 12'h000;
    rom[15488] = 12'h000;
    rom[15489] = 12'h000;
    rom[15490] = 12'h000;
    rom[15491] = 12'h000;
    rom[15492] = 12'h000;
    rom[15493] = 12'h000;
    rom[15494] = 12'h000;
    rom[15495] = 12'h000;
    rom[15496] = 12'h000;
    rom[15497] = 12'h000;
    rom[15498] = 12'h000;
    rom[15499] = 12'h000;
    rom[15500] = 12'h000;
    rom[15501] = 12'h000;
    rom[15502] = 12'h000;
    rom[15503] = 12'h000;
    rom[15504] = 12'h000;
    rom[15505] = 12'h000;
    rom[15506] = 12'h000;
    rom[15507] = 12'h000;
    rom[15508] = 12'h000;
    rom[15509] = 12'h000;
    rom[15510] = 12'h000;
    rom[15511] = 12'h000;
    rom[15512] = 12'h000;
    rom[15513] = 12'h000;
    rom[15514] = 12'h000;
    rom[15515] = 12'h000;
    rom[15516] = 12'h000;
    rom[15517] = 12'h000;
    rom[15518] = 12'h000;
    rom[15519] = 12'h000;
    rom[15520] = 12'h000;
    rom[15521] = 12'h000;
    rom[15522] = 12'h000;
    rom[15523] = 12'h000;
    rom[15524] = 12'h1ed;
    rom[15525] = 12'h1ed;
    rom[15526] = 12'h1ed;
    rom[15527] = 12'h1ed;
    rom[15528] = 12'h1ed;
    rom[15529] = 12'h2dd;
    rom[15530] = 12'h2dd;
    rom[15531] = 12'h2dd;
    rom[15532] = 12'h2dc;
    rom[15533] = 12'h2dc;
    rom[15534] = 12'h2dc;
    rom[15535] = 12'h2dc;
    rom[15536] = 12'h2dc;
    rom[15537] = 12'h2dc;
    rom[15538] = 12'h2dc;
    rom[15539] = 12'h2db;
    rom[15540] = 12'h2db;
    rom[15541] = 12'h2db;
    rom[15542] = 12'h2db;
    rom[15543] = 12'h3db;
    rom[15544] = 12'h3db;
    rom[15545] = 12'h3da;
    rom[15546] = 12'h3da;
    rom[15547] = 12'h3ca;
    rom[15548] = 12'h3ca;
    rom[15549] = 12'h3ca;
    rom[15550] = 12'h3ca;
    rom[15551] = 12'h3ca;
    rom[15552] = 12'h3ca;
    rom[15553] = 12'h3ca;
    rom[15554] = 12'h3ca;
    rom[15555] = 12'h3ca;
    rom[15556] = 12'h3c9;
    rom[15557] = 12'h3c9;
    rom[15558] = 12'h3c9;
    rom[15559] = 12'h3c9;
    rom[15560] = 12'h3c8;
    rom[15561] = 12'h3c8;
    rom[15562] = 12'h3c8;
    rom[15563] = 12'h3c8;
    rom[15564] = 12'h3c8;
    rom[15565] = 12'h3c7;
    rom[15566] = 12'h3b7;
    rom[15567] = 12'h3b7;
    rom[15568] = 12'h3b7;
    rom[15569] = 12'h3b6;
    rom[15570] = 12'h3b6;
    rom[15571] = 12'h3b6;
    rom[15572] = 12'h3b6;
    rom[15573] = 12'h3b5;
    rom[15574] = 12'h3b5;
    rom[15575] = 12'h3b5;
    rom[15576] = 12'h3b5;
    rom[15577] = 12'h3b5;
    rom[15578] = 12'h3a4;
    rom[15579] = 12'h3a4;
    rom[15580] = 12'h000;
    rom[15581] = 12'h000;
    rom[15582] = 12'h000;
    rom[15583] = 12'h000;
    rom[15584] = 12'h000;
    rom[15585] = 12'h000;
    rom[15586] = 12'h000;
    rom[15587] = 12'h000;
    rom[15588] = 12'h000;
    rom[15589] = 12'h000;
    rom[15590] = 12'h000;
    rom[15591] = 12'h000;
    rom[15592] = 12'h000;
    rom[15593] = 12'h000;
    rom[15594] = 12'h000;
    rom[15595] = 12'h000;
    rom[15596] = 12'h000;
    rom[15597] = 12'h000;
    rom[15598] = 12'h000;
    rom[15599] = 12'h000;
    rom[15600] = 12'h000;
    rom[15601] = 12'h000;
    rom[15602] = 12'h000;
    rom[15603] = 12'h000;
    rom[15604] = 12'h000;
    rom[15605] = 12'h000;
    rom[15606] = 12'h000;
    rom[15607] = 12'h000;
    rom[15608] = 12'h000;
    rom[15609] = 12'h000;
    rom[15610] = 12'h000;
    rom[15611] = 12'h000;
    rom[15612] = 12'h000;
    rom[15613] = 12'h000;
    rom[15614] = 12'h000;
    rom[15615] = 12'h000;
    rom[15616] = 12'h000;
    rom[15617] = 12'h000;
    rom[15618] = 12'h000;
    rom[15619] = 12'h000;
    rom[15620] = 12'h000;
    rom[15621] = 12'h000;
    rom[15622] = 12'h000;
    rom[15623] = 12'h000;
    rom[15624] = 12'h000;
    rom[15625] = 12'h000;
    rom[15626] = 12'h000;
    rom[15627] = 12'h000;
    rom[15628] = 12'h000;
    rom[15629] = 12'h000;
    rom[15630] = 12'h000;
    rom[15631] = 12'h000;
    rom[15632] = 12'h000;
    rom[15633] = 12'h000;
    rom[15634] = 12'h000;
    rom[15635] = 12'h000;
    rom[15636] = 12'h000;
    rom[15637] = 12'h000;
    rom[15638] = 12'h000;
    rom[15639] = 12'h000;
    rom[15640] = 12'h000;
    rom[15641] = 12'h000;
    rom[15642] = 12'h000;
    rom[15643] = 12'h000;
    rom[15644] = 12'h000;
    rom[15645] = 12'h000;
    rom[15646] = 12'h000;
    rom[15647] = 12'h000;
    rom[15648] = 12'h000;
    rom[15649] = 12'h000;
    rom[15650] = 12'h000;
    rom[15651] = 12'h000;
    rom[15652] = 12'h000;
    rom[15653] = 12'h000;
    rom[15654] = 12'h1ed;
    rom[15655] = 12'h1ed;
    rom[15656] = 12'h2ed;
    rom[15657] = 12'h2dd;
    rom[15658] = 12'h2dd;
    rom[15659] = 12'h2dd;
    rom[15660] = 12'h2dc;
    rom[15661] = 12'h2dc;
    rom[15662] = 12'h2dc;
    rom[15663] = 12'h2dc;
    rom[15664] = 12'h2dc;
    rom[15665] = 12'h2dc;
    rom[15666] = 12'h2dc;
    rom[15667] = 12'h2db;
    rom[15668] = 12'h2db;
    rom[15669] = 12'h2db;
    rom[15670] = 12'h3db;
    rom[15671] = 12'h3db;
    rom[15672] = 12'h3da;
    rom[15673] = 12'h3da;
    rom[15674] = 12'h3da;
    rom[15675] = 12'h3ca;
    rom[15676] = 12'h3ca;
    rom[15677] = 12'h3ca;
    rom[15678] = 12'h3ca;
    rom[15679] = 12'h3ca;
    rom[15680] = 12'h3ca;
    rom[15681] = 12'h3ca;
    rom[15682] = 12'h3ca;
    rom[15683] = 12'h3ca;
    rom[15684] = 12'h3c9;
    rom[15685] = 12'h3c9;
    rom[15686] = 12'h3c9;
    rom[15687] = 12'h3c9;
    rom[15688] = 12'h3c8;
    rom[15689] = 12'h3c8;
    rom[15690] = 12'h3c8;
    rom[15691] = 12'h3c8;
    rom[15692] = 12'h3c8;
    rom[15693] = 12'h3c7;
    rom[15694] = 12'h3b7;
    rom[15695] = 12'h3b7;
    rom[15696] = 12'h3b7;
    rom[15697] = 12'h3b6;
    rom[15698] = 12'h3b6;
    rom[15699] = 12'h3b6;
    rom[15700] = 12'h3b6;
    rom[15701] = 12'h3b6;
    rom[15702] = 12'h3b5;
    rom[15703] = 12'h3b5;
    rom[15704] = 12'h3b5;
    rom[15705] = 12'h3b5;
    rom[15706] = 12'h000;
    rom[15707] = 12'h000;
    rom[15708] = 12'h000;
    rom[15709] = 12'h000;
    rom[15710] = 12'h000;
    rom[15711] = 12'h000;
    rom[15712] = 12'h000;
    rom[15713] = 12'h000;
    rom[15714] = 12'h000;
    rom[15715] = 12'h000;
    rom[15716] = 12'h000;
    rom[15717] = 12'h000;
    rom[15718] = 12'h000;
    rom[15719] = 12'h000;
    rom[15720] = 12'h000;
    rom[15721] = 12'h000;
    rom[15722] = 12'h000;
    rom[15723] = 12'h000;
    rom[15724] = 12'h000;
    rom[15725] = 12'h000;
    rom[15726] = 12'h000;
    rom[15727] = 12'h000;
    rom[15728] = 12'h000;
    rom[15729] = 12'h000;
    rom[15730] = 12'h000;
    rom[15731] = 12'h000;
    rom[15732] = 12'h000;
    rom[15733] = 12'h000;
    rom[15734] = 12'h000;
    rom[15735] = 12'h000;
    rom[15736] = 12'h000;
    rom[15737] = 12'h000;
    rom[15738] = 12'h000;
    rom[15739] = 12'h000;
    rom[15740] = 12'h000;
    rom[15741] = 12'h000;
    rom[15742] = 12'h000;
    rom[15743] = 12'h000;
    rom[15744] = 12'h000;
    rom[15745] = 12'h000;
    rom[15746] = 12'h000;
    rom[15747] = 12'h000;
    rom[15748] = 12'h000;
    rom[15749] = 12'h000;
    rom[15750] = 12'h000;
    rom[15751] = 12'h000;
    rom[15752] = 12'h000;
    rom[15753] = 12'h000;
    rom[15754] = 12'h000;
    rom[15755] = 12'h000;
    rom[15756] = 12'h000;
    rom[15757] = 12'h000;
    rom[15758] = 12'h000;
    rom[15759] = 12'h000;
    rom[15760] = 12'h000;
    rom[15761] = 12'h000;
    rom[15762] = 12'h000;
    rom[15763] = 12'h000;
    rom[15764] = 12'h000;
    rom[15765] = 12'h000;
    rom[15766] = 12'h000;
    rom[15767] = 12'h000;
    rom[15768] = 12'h000;
    rom[15769] = 12'h000;
    rom[15770] = 12'h000;
    rom[15771] = 12'h000;
    rom[15772] = 12'h000;
    rom[15773] = 12'h000;
    rom[15774] = 12'h000;
    rom[15775] = 12'h000;
    rom[15776] = 12'h000;
    rom[15777] = 12'h000;
    rom[15778] = 12'h000;
    rom[15779] = 12'h000;
    rom[15780] = 12'h000;
    rom[15781] = 12'h000;
    rom[15782] = 12'h000;
    rom[15783] = 12'h000;
    rom[15784] = 12'h1ed;
    rom[15785] = 12'h2dd;
    rom[15786] = 12'h2dd;
    rom[15787] = 12'h2dd;
    rom[15788] = 12'h2dc;
    rom[15789] = 12'h2dc;
    rom[15790] = 12'h2dc;
    rom[15791] = 12'h2dc;
    rom[15792] = 12'h2dc;
    rom[15793] = 12'h2dc;
    rom[15794] = 12'h2db;
    rom[15795] = 12'h2db;
    rom[15796] = 12'h2db;
    rom[15797] = 12'h2db;
    rom[15798] = 12'h3db;
    rom[15799] = 12'h3db;
    rom[15800] = 12'h3da;
    rom[15801] = 12'h3da;
    rom[15802] = 12'h3ca;
    rom[15803] = 12'h3ca;
    rom[15804] = 12'h3ca;
    rom[15805] = 12'h3ca;
    rom[15806] = 12'h3ca;
    rom[15807] = 12'h3ca;
    rom[15808] = 12'h3ca;
    rom[15809] = 12'h3ca;
    rom[15810] = 12'h3ca;
    rom[15811] = 12'h3ca;
    rom[15812] = 12'h3c9;
    rom[15813] = 12'h3c9;
    rom[15814] = 12'h3c9;
    rom[15815] = 12'h3c9;
    rom[15816] = 12'h3c9;
    rom[15817] = 12'h3c8;
    rom[15818] = 12'h3c8;
    rom[15819] = 12'h3c8;
    rom[15820] = 12'h3c8;
    rom[15821] = 12'h3c7;
    rom[15822] = 12'h3b7;
    rom[15823] = 12'h3b7;
    rom[15824] = 12'h3b7;
    rom[15825] = 12'h3b7;
    rom[15826] = 12'h3b6;
    rom[15827] = 12'h3b6;
    rom[15828] = 12'h3b6;
    rom[15829] = 12'h3b6;
    rom[15830] = 12'h3b5;
    rom[15831] = 12'h000;
    rom[15832] = 12'h000;
    rom[15833] = 12'h000;
    rom[15834] = 12'h000;
    rom[15835] = 12'h000;
    rom[15836] = 12'h000;
    rom[15837] = 12'h000;
    rom[15838] = 12'h000;
    rom[15839] = 12'h000;
    rom[15840] = 12'h000;
    rom[15841] = 12'h000;
    rom[15842] = 12'h000;
    rom[15843] = 12'h000;
    rom[15844] = 12'h000;
    rom[15845] = 12'h000;
    rom[15846] = 12'h000;
    rom[15847] = 12'h000;
    rom[15848] = 12'h000;
    rom[15849] = 12'h000;
    rom[15850] = 12'h000;
    rom[15851] = 12'h000;
    rom[15852] = 12'h000;
    rom[15853] = 12'h000;
    rom[15854] = 12'h000;
    rom[15855] = 12'h000;
    rom[15856] = 12'h000;
    rom[15857] = 12'h000;
    rom[15858] = 12'h000;
    rom[15859] = 12'h000;
    rom[15860] = 12'h000;
    rom[15861] = 12'h000;
    rom[15862] = 12'h000;
    rom[15863] = 12'h000;
    rom[15864] = 12'h000;
    rom[15865] = 12'h000;
    rom[15866] = 12'h000;
    rom[15867] = 12'h000;
    rom[15868] = 12'h000;
    rom[15869] = 12'h000;
    rom[15870] = 12'h000;
    rom[15871] = 12'h000;
    rom[15872] = 12'h000;
    rom[15873] = 12'h000;
    rom[15874] = 12'h000;
    rom[15875] = 12'h000;
    rom[15876] = 12'h000;
    rom[15877] = 12'h000;
    rom[15878] = 12'h000;
    rom[15879] = 12'h000;
    rom[15880] = 12'h000;
    rom[15881] = 12'h000;
    rom[15882] = 12'h000;
    rom[15883] = 12'h000;
    rom[15884] = 12'h000;
    rom[15885] = 12'h000;
    rom[15886] = 12'h000;
    rom[15887] = 12'h000;
    rom[15888] = 12'h000;
    rom[15889] = 12'h000;
    rom[15890] = 12'h000;
    rom[15891] = 12'h000;
    rom[15892] = 12'h000;
    rom[15893] = 12'h000;
    rom[15894] = 12'h000;
    rom[15895] = 12'h000;
    rom[15896] = 12'h000;
    rom[15897] = 12'h000;
    rom[15898] = 12'h000;
    rom[15899] = 12'h000;
    rom[15900] = 12'h000;
    rom[15901] = 12'h000;
    rom[15902] = 12'h000;
    rom[15903] = 12'h000;
    rom[15904] = 12'h000;
    rom[15905] = 12'h000;
    rom[15906] = 12'h000;
    rom[15907] = 12'h000;
    rom[15908] = 12'h000;
    rom[15909] = 12'h000;
    rom[15910] = 12'h000;
    rom[15911] = 12'h000;
    rom[15912] = 12'h000;
    rom[15913] = 12'h000;
    rom[15914] = 12'h000;
    rom[15915] = 12'h2dc;
    rom[15916] = 12'h2dc;
    rom[15917] = 12'h2dc;
    rom[15918] = 12'h2dc;
    rom[15919] = 12'h2dc;
    rom[15920] = 12'h2dc;
    rom[15921] = 12'h2dc;
    rom[15922] = 12'h2db;
    rom[15923] = 12'h2db;
    rom[15924] = 12'h2db;
    rom[15925] = 12'h2db;
    rom[15926] = 12'h3db;
    rom[15927] = 12'h3db;
    rom[15928] = 12'h3da;
    rom[15929] = 12'h3da;
    rom[15930] = 12'h3ca;
    rom[15931] = 12'h3ca;
    rom[15932] = 12'h3ca;
    rom[15933] = 12'h3ca;
    rom[15934] = 12'h3ca;
    rom[15935] = 12'h3ca;
    rom[15936] = 12'h3ca;
    rom[15937] = 12'h3ca;
    rom[15938] = 12'h3ca;
    rom[15939] = 12'h3ca;
    rom[15940] = 12'h3ca;
    rom[15941] = 12'h3c9;
    rom[15942] = 12'h3c9;
    rom[15943] = 12'h3c9;
    rom[15944] = 12'h3c9;
    rom[15945] = 12'h3c8;
    rom[15946] = 12'h3c8;
    rom[15947] = 12'h3c8;
    rom[15948] = 12'h3c8;
    rom[15949] = 12'h3c7;
    rom[15950] = 12'h3b7;
    rom[15951] = 12'h3b7;
    rom[15952] = 12'h3b7;
    rom[15953] = 12'h3b7;
    rom[15954] = 12'h3b6;
    rom[15955] = 12'h3b6;
    rom[15956] = 12'h3b6;
    rom[15957] = 12'h000;
    rom[15958] = 12'h000;
    rom[15959] = 12'h000;
    rom[15960] = 12'h000;
    rom[15961] = 12'h000;
    rom[15962] = 12'h000;
    rom[15963] = 12'h000;
    rom[15964] = 12'h000;
    rom[15965] = 12'h000;
    rom[15966] = 12'h000;
    rom[15967] = 12'h000;
    rom[15968] = 12'h000;
    rom[15969] = 12'h000;
    rom[15970] = 12'h000;
    rom[15971] = 12'h000;
    rom[15972] = 12'h000;
    rom[15973] = 12'h000;
    rom[15974] = 12'h000;
    rom[15975] = 12'h000;
    rom[15976] = 12'h000;
    rom[15977] = 12'h000;
    rom[15978] = 12'h000;
    rom[15979] = 12'h000;
    rom[15980] = 12'h000;
    rom[15981] = 12'h000;
    rom[15982] = 12'h000;
    rom[15983] = 12'h000;
    rom[15984] = 12'h000;
    rom[15985] = 12'h000;
    rom[15986] = 12'h000;
    rom[15987] = 12'h000;
    rom[15988] = 12'h000;
    rom[15989] = 12'h000;
    rom[15990] = 12'h000;
    rom[15991] = 12'h000;
    rom[15992] = 12'h000;
    rom[15993] = 12'h000;
    rom[15994] = 12'h000;
    rom[15995] = 12'h000;
    rom[15996] = 12'h000;
    rom[15997] = 12'h000;
    rom[15998] = 12'h000;
    rom[15999] = 12'h000;
    rom[16000] = 12'h000;
    rom[16001] = 12'h000;
    rom[16002] = 12'h000;
    rom[16003] = 12'h000;
    rom[16004] = 12'h000;
    rom[16005] = 12'h000;
    rom[16006] = 12'h000;
    rom[16007] = 12'h000;
    rom[16008] = 12'h000;
    rom[16009] = 12'h000;
    rom[16010] = 12'h000;
    rom[16011] = 12'h000;
    rom[16012] = 12'h000;
    rom[16013] = 12'h000;
    rom[16014] = 12'h000;
    rom[16015] = 12'h000;
    rom[16016] = 12'h000;
    rom[16017] = 12'h000;
    rom[16018] = 12'h000;
    rom[16019] = 12'h000;
    rom[16020] = 12'h000;
    rom[16021] = 12'h000;
    rom[16022] = 12'h000;
    rom[16023] = 12'h000;
    rom[16024] = 12'h000;
    rom[16025] = 12'h000;
    rom[16026] = 12'h000;
    rom[16027] = 12'h000;
    rom[16028] = 12'h000;
    rom[16029] = 12'h000;
    rom[16030] = 12'h000;
    rom[16031] = 12'h000;
    rom[16032] = 12'h000;
    rom[16033] = 12'h000;
    rom[16034] = 12'h000;
    rom[16035] = 12'h000;
    rom[16036] = 12'h000;
    rom[16037] = 12'h000;
    rom[16038] = 12'h000;
    rom[16039] = 12'h000;
    rom[16040] = 12'h000;
    rom[16041] = 12'h000;
    rom[16042] = 12'h000;
    rom[16043] = 12'h000;
    rom[16044] = 12'h000;
    rom[16045] = 12'h000;
    rom[16046] = 12'h2dc;
    rom[16047] = 12'h2dc;
    rom[16048] = 12'h2dc;
    rom[16049] = 12'h2db;
    rom[16050] = 12'h2db;
    rom[16051] = 12'h2db;
    rom[16052] = 12'h2db;
    rom[16053] = 12'h3db;
    rom[16054] = 12'h3db;
    rom[16055] = 12'h3da;
    rom[16056] = 12'h3da;
    rom[16057] = 12'h3ca;
    rom[16058] = 12'h3ca;
    rom[16059] = 12'h3ca;
    rom[16060] = 12'h3ca;
    rom[16061] = 12'h3ca;
    rom[16062] = 12'h3ca;
    rom[16063] = 12'h3ca;
    rom[16064] = 12'h3ca;
    rom[16065] = 12'h3ca;
    rom[16066] = 12'h3ca;
    rom[16067] = 12'h3ca;
    rom[16068] = 12'h3ca;
    rom[16069] = 12'h3c9;
    rom[16070] = 12'h3c9;
    rom[16071] = 12'h3c9;
    rom[16072] = 12'h3c9;
    rom[16073] = 12'h3c8;
    rom[16074] = 12'h3c8;
    rom[16075] = 12'h3c8;
    rom[16076] = 12'h3c8;
    rom[16077] = 12'h3c7;
    rom[16078] = 12'h3b7;
    rom[16079] = 12'h3b7;
    rom[16080] = 12'h3b7;
    rom[16081] = 12'h3b7;
    rom[16082] = 12'h000;
    rom[16083] = 12'h000;
    rom[16084] = 12'h000;
    rom[16085] = 12'h000;
    rom[16086] = 12'h000;
    rom[16087] = 12'h000;
    rom[16088] = 12'h000;
    rom[16089] = 12'h000;
    rom[16090] = 12'h000;
    rom[16091] = 12'h000;
    rom[16092] = 12'h000;
    rom[16093] = 12'h000;
    rom[16094] = 12'h000;
    rom[16095] = 12'h000;
    rom[16096] = 12'h000;
    rom[16097] = 12'h000;
    rom[16098] = 12'h000;
    rom[16099] = 12'h000;
    rom[16100] = 12'h000;
    rom[16101] = 12'h000;
    rom[16102] = 12'h000;
    rom[16103] = 12'h000;
    rom[16104] = 12'h000;
    rom[16105] = 12'h000;
    rom[16106] = 12'h000;
    rom[16107] = 12'h000;
    rom[16108] = 12'h000;
    rom[16109] = 12'h000;
    rom[16110] = 12'h000;
    rom[16111] = 12'h000;
    rom[16112] = 12'h000;
    rom[16113] = 12'h000;
    rom[16114] = 12'h000;
    rom[16115] = 12'h000;
    rom[16116] = 12'h000;
    rom[16117] = 12'h000;
    rom[16118] = 12'h000;
    rom[16119] = 12'h000;
    rom[16120] = 12'h000;
    rom[16121] = 12'h000;
    rom[16122] = 12'h000;
    rom[16123] = 12'h000;
    rom[16124] = 12'h000;
    rom[16125] = 12'h000;
    rom[16126] = 12'h000;
    rom[16127] = 12'h000;
    rom[16128] = 12'h000;
    rom[16129] = 12'h000;
    rom[16130] = 12'h000;
    rom[16131] = 12'h000;
    rom[16132] = 12'h000;
    rom[16133] = 12'h000;
    rom[16134] = 12'h000;
    rom[16135] = 12'h000;
    rom[16136] = 12'h000;
    rom[16137] = 12'h000;
    rom[16138] = 12'h000;
    rom[16139] = 12'h000;
    rom[16140] = 12'h000;
    rom[16141] = 12'h000;
    rom[16142] = 12'h000;
    rom[16143] = 12'h000;
    rom[16144] = 12'h000;
    rom[16145] = 12'h000;
    rom[16146] = 12'h000;
    rom[16147] = 12'h000;
    rom[16148] = 12'h000;
    rom[16149] = 12'h000;
    rom[16150] = 12'h000;
    rom[16151] = 12'h000;
    rom[16152] = 12'h000;
    rom[16153] = 12'h000;
    rom[16154] = 12'h000;
    rom[16155] = 12'h000;
    rom[16156] = 12'h000;
    rom[16157] = 12'h000;
    rom[16158] = 12'h000;
    rom[16159] = 12'h000;
    rom[16160] = 12'h000;
    rom[16161] = 12'h000;
    rom[16162] = 12'h000;
    rom[16163] = 12'h000;
    rom[16164] = 12'h000;
    rom[16165] = 12'h000;
    rom[16166] = 12'h000;
    rom[16167] = 12'h000;
    rom[16168] = 12'h000;
    rom[16169] = 12'h000;
    rom[16170] = 12'h000;
    rom[16171] = 12'h000;
    rom[16172] = 12'h000;
    rom[16173] = 12'h000;
    rom[16174] = 12'h000;
    rom[16175] = 12'h000;
    rom[16176] = 12'h000;
    rom[16177] = 12'h000;
    rom[16178] = 12'h2db;
    rom[16179] = 12'h2db;
    rom[16180] = 12'h2db;
    rom[16181] = 12'h3db;
    rom[16182] = 12'h3db;
    rom[16183] = 12'h3da;
    rom[16184] = 12'h3da;
    rom[16185] = 12'h3ca;
    rom[16186] = 12'h3ca;
    rom[16187] = 12'h3ca;
    rom[16188] = 12'h3ca;
    rom[16189] = 12'h3ca;
    rom[16190] = 12'h3ca;
    rom[16191] = 12'h3ca;
    rom[16192] = 12'h3ca;
    rom[16193] = 12'h3ca;
    rom[16194] = 12'h3ca;
    rom[16195] = 12'h3ca;
    rom[16196] = 12'h3ca;
    rom[16197] = 12'h3c9;
    rom[16198] = 12'h3c9;
    rom[16199] = 12'h3c9;
    rom[16200] = 12'h3c9;
    rom[16201] = 12'h3c8;
    rom[16202] = 12'h3c8;
    rom[16203] = 12'h3c8;
    rom[16204] = 12'h3c8;
    rom[16205] = 12'h4b8;
    rom[16206] = 12'h000;
    rom[16207] = 12'h000;
    rom[16208] = 12'h000;
    rom[16209] = 12'h000;
    rom[16210] = 12'h000;
    rom[16211] = 12'h000;
    rom[16212] = 12'h000;
    rom[16213] = 12'h000;
    rom[16214] = 12'h000;
    rom[16215] = 12'h000;
    rom[16216] = 12'h000;
    rom[16217] = 12'h000;
    rom[16218] = 12'h000;
    rom[16219] = 12'h000;
    rom[16220] = 12'h000;
    rom[16221] = 12'h000;
    rom[16222] = 12'h000;
    rom[16223] = 12'h000;
    rom[16224] = 12'h000;
    rom[16225] = 12'h000;
    rom[16226] = 12'h000;
    rom[16227] = 12'h000;
    rom[16228] = 12'h000;
    rom[16229] = 12'h000;
    rom[16230] = 12'h000;
    rom[16231] = 12'h000;
    rom[16232] = 12'h000;
    rom[16233] = 12'h000;
    rom[16234] = 12'h000;
    rom[16235] = 12'h000;
    rom[16236] = 12'h000;
    rom[16237] = 12'h000;
    rom[16238] = 12'h000;
    rom[16239] = 12'h000;
    rom[16240] = 12'h000;
    rom[16241] = 12'h000;
    rom[16242] = 12'h000;
    rom[16243] = 12'h000;
    rom[16244] = 12'h000;
    rom[16245] = 12'h000;
    rom[16246] = 12'h000;
    rom[16247] = 12'h000;
    rom[16248] = 12'h000;
    rom[16249] = 12'h000;
    rom[16250] = 12'h000;
    rom[16251] = 12'h000;
    rom[16252] = 12'h000;
    rom[16253] = 12'h000;
    rom[16254] = 12'h000;
    rom[16255] = 12'h000;
    rom[16256] = 12'h000;
    rom[16257] = 12'h000;
    rom[16258] = 12'h000;
    rom[16259] = 12'h000;
    rom[16260] = 12'h000;
    rom[16261] = 12'h000;
    rom[16262] = 12'h000;
    rom[16263] = 12'h000;
    rom[16264] = 12'h000;
    rom[16265] = 12'h000;
    rom[16266] = 12'h000;
    rom[16267] = 12'h000;
    rom[16268] = 12'h000;
    rom[16269] = 12'h000;
    rom[16270] = 12'h000;
    rom[16271] = 12'h000;
    rom[16272] = 12'h000;
    rom[16273] = 12'h000;
    rom[16274] = 12'h000;
    rom[16275] = 12'h000;
    rom[16276] = 12'h000;
    rom[16277] = 12'h000;
    rom[16278] = 12'h000;
    rom[16279] = 12'h000;
    rom[16280] = 12'h000;
    rom[16281] = 12'h000;
    rom[16282] = 12'h000;
    rom[16283] = 12'h000;
    rom[16284] = 12'h000;
    rom[16285] = 12'h000;
    rom[16286] = 12'h000;
    rom[16287] = 12'h000;
    rom[16288] = 12'h000;
    rom[16289] = 12'h000;
    rom[16290] = 12'h000;
    rom[16291] = 12'h000;
    rom[16292] = 12'h000;
    rom[16293] = 12'h000;
    rom[16294] = 12'h000;
    rom[16295] = 12'h000;
    rom[16296] = 12'h000;
    rom[16297] = 12'h000;
    rom[16298] = 12'h000;
    rom[16299] = 12'h000;
    rom[16300] = 12'h000;
    rom[16301] = 12'h000;
    rom[16302] = 12'h000;
    rom[16303] = 12'h000;
    rom[16304] = 12'h000;
    rom[16305] = 12'h000;
    rom[16306] = 12'h000;
    rom[16307] = 12'h000;
    rom[16308] = 12'h000;
    rom[16309] = 12'h000;
    rom[16310] = 12'h000;
    rom[16311] = 12'h0f0;
    rom[16312] = 12'h3da;
    rom[16313] = 12'h3ca;
    rom[16314] = 12'h3ca;
    rom[16315] = 12'h3ca;
    rom[16316] = 12'h3ca;
    rom[16317] = 12'h3ca;
    rom[16318] = 12'h3ca;
    rom[16319] = 12'h3ca;
    rom[16320] = 12'h3ca;
    rom[16321] = 12'h3ca;
    rom[16322] = 12'h3ca;
    rom[16323] = 12'h3ca;
    rom[16324] = 12'h3ca;
    rom[16325] = 12'h3c9;
    rom[16326] = 12'h3c9;
    rom[16327] = 12'h3c9;
    rom[16328] = 12'h000;
    rom[16329] = 12'h000;
    rom[16330] = 12'h000;
    rom[16331] = 12'h000;
    rom[16332] = 12'h000;
    rom[16333] = 12'h000;
    rom[16334] = 12'h000;
    rom[16335] = 12'h000;
    rom[16336] = 12'h000;
    rom[16337] = 12'h000;
    rom[16338] = 12'h000;
    rom[16339] = 12'h000;
    rom[16340] = 12'h000;
    rom[16341] = 12'h000;
    rom[16342] = 12'h000;
    rom[16343] = 12'h000;
    rom[16344] = 12'h000;
    rom[16345] = 12'h000;
    rom[16346] = 12'h000;
    rom[16347] = 12'h000;
    rom[16348] = 12'h000;
    rom[16349] = 12'h000;
    rom[16350] = 12'h000;
    rom[16351] = 12'h000;
    rom[16352] = 12'h000;
    rom[16353] = 12'h000;
    rom[16354] = 12'h000;
    rom[16355] = 12'h000;
    rom[16356] = 12'h000;
    rom[16357] = 12'h000;
    rom[16358] = 12'h000;
    rom[16359] = 12'h000;
    rom[16360] = 12'h000;
    rom[16361] = 12'h000;
    rom[16362] = 12'h000;
    rom[16363] = 12'h000;
    rom[16364] = 12'h000;
    rom[16365] = 12'h000;
    rom[16366] = 12'h000;
    rom[16367] = 12'h000;
    rom[16368] = 12'h000;
    rom[16369] = 12'h000;
    rom[16370] = 12'h000;
    rom[16371] = 12'h000;
    rom[16372] = 12'h000;
    rom[16373] = 12'h000;
    rom[16374] = 12'h000;
    rom[16375] = 12'h000;
    rom[16376] = 12'h000;
    rom[16377] = 12'h000;
    rom[16378] = 12'h000;
    rom[16379] = 12'h000;
    rom[16380] = 12'h000;
    rom[16381] = 12'h000;
    rom[16382] = 12'h000;
    rom[16383] = 12'h000;
    */
  end

endmodule